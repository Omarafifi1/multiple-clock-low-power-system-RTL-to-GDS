module DLY3X1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module DLY2X1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module DLY4X1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX40M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX5M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVXLM (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX32M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX40M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX16M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module TIEHIM (
	Y, 
	VDD, 
	VSS);
   output Y;
   inout VDD;
   inout VSS;
endmodule

module TIELOM (
	Y, 
	VDD, 
	VSS);
   output Y;
   inout VDD;
   inout VSS;
endmodule

module CLKAND2X12M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI21BX4M (
	Y, 
	B0N, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0N;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKNAND2X4M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2X3M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2X4M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND3X3M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB1X2M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module NAND4X2M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKAND2X6M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2X3M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKNAND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module XNOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2BX4M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AND2X4M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI2B1X2M (
	Y, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module MXI2X1M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB2X1M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module AND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MXI2X2M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI2B1X4M (
	Y, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module XOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2B1X4M (
	Y, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI21X4M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI2B1X2M (
	Y, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module CLKNAND2X8M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2BX8M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module MXI2X6M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND3X4M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MXI2X4M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2X4M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND3BX4M (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NOR2BX8M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AND2X12M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2X6M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module XNOR2X4M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI211X4M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND2X5M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AO21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI21X1M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR2BX2M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NAND2BX2M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module OAI2B11X4M (
	Y, 
	C0, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module XOR2X4M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI2B1X8M (
	Y, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module MX2X2M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2X8M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI22X1M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI22X1M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI2B1X8M (
	Y, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR2X8M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI2BB1X4M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module XOR2X8M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2X6M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND3X1M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AO2B2X4M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module INVX3M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI21X4M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR3X4M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2X5M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKAND2X8M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND4X6M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND4X4M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND4X4M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB2X8M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module AND3X6M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND2X8M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2X12M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX8M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX10M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX8M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX10M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX8M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX6M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module SDFFRQX2M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFRX1M (
	SI, 
	SE, 
	RN, 
	QN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output QN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module NAND4BX1M (
	Y, 
	D, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NOR3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR4X1M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI211X2M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module DLY1X4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AO2B2X2M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI31X1M (
	Y, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI32X1M (
	Y, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AND3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI31X2M (
	Y, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI2BB2XLM (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module AOI33X2M (
	Y, 
	B2, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B2;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OA21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI222X1M (
	Y, 
	C1, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C1;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AO21XLM (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AO22X1M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module ADDHX1M (
	S, 
	CO, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB1X1M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module OR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module XNOR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR3X1M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI21X1M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND2BX1M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module CLKXOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2BX1M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module OAI2B2X1M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND4BBX1M (
	Y, 
	D, 
	C, 
	BN, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input BN;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module OR3X1M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI32X1M (
	Y, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AND2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND4X1M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR4XLM (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI33XLM (
	Y, 
	B2, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B2;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR3BX2M (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module XOR3XLM (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX12M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module SDFFRHQX4M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFRHQX2M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFSQX2M (
	SN, 
	SI, 
	SE, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SN;
   input SI;
   input SE;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFSQX1M (
	SN, 
	SI, 
	SE, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SN;
   input SI;
   input SE;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module AND3XLM (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX4XLM (
	Y, 
	S1, 
	S0, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S1;
   input S0;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX4X1M (
	Y, 
	S1, 
	S0, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S1;
   input S0;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module SDFFRQX4M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFRHQX1M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFRQX1M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module AND4X2M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND3BX2M (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AOI211X2M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI222X1M (
	Y, 
	C1, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C1;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI221XLM (
	Y, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI221X1M (
	Y, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI33X1M (
	Y, 
	B2, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B2;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI222X4M (
	Y, 
	C1, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C1;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI2B11X2M (
	Y, 
	C0, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI211X1M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI211X1M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OA21X1M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI31X1M (
	Y, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI2B11X1M (
	Y, 
	C0, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI2B1X1M (
	Y, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module ADDFHX2M (
	S, 
	CO, 
	CI, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input CI;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module ADDFX1M (
	S, 
	CO, 
	CI, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input CI;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module ADDFHX1M (
	S, 
	CO, 
	CI, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input CI;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX12M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKMX2X2M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2X6M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2X8M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module ADDFX2M (
	S, 
	CO, 
	CI, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input CI;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI21BX2M (
	Y, 
	B0N, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0N;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI21BX1M (
	Y, 
	B0N, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0N;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI2BB1X1M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module TLATNCAX3M (
	ECK, 
	E, 
	CK, 
	VDD, 
	VSS);
   output ECK;
   input E;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module NOR4BX1M (
	Y, 
	D, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Expert(TM) in wire load mode
// Version   : K-2015.06
// Date      : Thu Aug 29 00:22:05 2024
/////////////////////////////////////////////////////////////
module mux_2x1_0 (
	in0, 
	in1, 
	sel, 
	out, 
	VDD, 
	VSS);
   input in0;
   input in1;
   input sel;
   output out;
   inout VDD;
   inout VSS;

   // Module instantiations
   AO2B2X2M U1 (
	.Y(out),
	.B1(in1),
	.B0(sel),
	.A1N(sel),
	.A0(in0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux_2x1_6 (
	in0, 
	in1, 
	sel, 
	out, 
	VDD, 
	VSS);
   input in0;
   input in1;
   input sel;
   output out;
   inout VDD;
   inout VSS;

   // Module instantiations
   AO2B2X4M U1 (
	.Y(out),
	.B1(in1),
	.B0(sel),
	.A1N(sel),
	.A0(in0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux_2x1_5 (
	in0, 
	in1, 
	sel, 
	out, 
	VDD, 
	VSS);
   input in0;
   input in1;
   input sel;
   output out;
   inout VDD;
   inout VSS;

   // Module instantiations
   AO2B2X2M U1 (
	.Y(out),
	.B1(in1),
	.B0(sel),
	.A1N(sel),
	.A0(in0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux_2x1_4 (
	in0, 
	in1, 
	sel, 
	out, 
	VDD, 
	VSS);
   input in0;
   input in1;
   input sel;
   output out;
   inout VDD;
   inout VSS;

   // Module instantiations
   AO2B2X2M U1 (
	.Y(out),
	.B1(in1),
	.B0(sel),
	.A1N(sel),
	.A0(in0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux_2x1_3 (
	in0, 
	in1, 
	sel, 
	out, 
	VDD, 
	VSS);
   input in0;
   input in1;
   input sel;
   output out;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN6_rst_n;
   wire FE_PHN5_rst_n;
   wire FE_PHN3_SCAN_RST;
   wire FE_PHN0_SCAN_RST;

   // Module instantiations
   DLY4X1M FE_PHC6_rst_n (
	.Y(FE_PHN6_rst_n),
	.A(FE_PHN5_rst_n), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC5_rst_n (
	.Y(FE_PHN5_rst_n),
	.A(in0), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC3_SCAN_RST (
	.Y(FE_PHN3_SCAN_RST),
	.A(FE_PHN0_SCAN_RST), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC0_SCAN_RST (
	.Y(FE_PHN0_SCAN_RST),
	.A(in1), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U1 (
	.Y(out),
	.B1(FE_PHN3_SCAN_RST),
	.B0(sel),
	.A1N(sel),
	.A0(FE_PHN6_rst_n), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux_2x1_2 (
	in0, 
	in1, 
	sel, 
	out, 
	VDD, 
	VSS);
   input in0;
   input in1;
   input sel;
   output out;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN4_SCAN_RST;
   wire FE_PHN2_SCAN_RST;

   // Module instantiations
   DLY4X1M FE_PHC4_SCAN_RST (
	.Y(FE_PHN4_SCAN_RST),
	.A(FE_PHN2_SCAN_RST), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC2_SCAN_RST (
	.Y(FE_PHN2_SCAN_RST),
	.A(in1), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U1 (
	.Y(out),
	.B1(FE_PHN4_SCAN_RST),
	.B0(sel),
	.A1N(sel),
	.A0(in0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux_2x1_1 (
	in0, 
	in1, 
	sel, 
	out, 
	VDD, 
	VSS);
   input in0;
   input in1;
   input sel;
   output out;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN1_SCAN_RST;

   // Module instantiations
   DLY4X1M FE_PHC1_SCAN_RST (
	.Y(FE_PHN1_SCAN_RST),
	.A(in1), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U1 (
	.Y(out),
	.B1(FE_PHN1_SCAN_RST),
	.B0(sel),
	.A1N(sel),
	.A0(in0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module sys_ctrl_test_1 (
	clk, 
	rst_n, 
	alu_out, 
	out_valid, 
	rx_P_data, 
	rx_d_valid, 
	full_flag, 
	rd_data, 
	rd_data_valid, 
	alu_en, 
	alu_fun, 
	clk_en, 
	address, 
	w_en, 
	r_en, 
	w_data, 
	tx_P_data, 
	w_inc, 
	clk_div_en, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN2_scan_rst_sync1_mux_out, 
	VDD, 
	VSS);
   input clk;
   input rst_n;
   input [15:0] alu_out;
   input out_valid;
   input [7:0] rx_P_data;
   input rx_d_valid;
   input full_flag;
   input [7:0] rd_data;
   input rd_data_valid;
   output alu_en;
   output [3:0] alu_fun;
   output clk_en;
   output [3:0] address;
   output w_en;
   output r_en;
   output [7:0] w_data;
   output [7:0] tx_P_data;
   output w_inc;
   output clk_div_en;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN2_scan_rst_sync1_mux_out;
   inout VDD;
   inout VSS;

   // Internal wires
   wire LTIE_LTIELO_NET;
   wire FE_OFN12_address_3_;
   wire n17;
   wire n18;
   wire n19;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n15;
   wire n16;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire [3:0] current_state;

   assign test_so = n99 ;

   // Module instantiations
   TIELOM LTIE_LTIELO (
	.Y(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M FE_OFC12_address_3_ (
	.Y(address[3]),
	.A(FE_OFN12_address_3_), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \address_reg[1]  (
	.SI(n19),
	.SE(test_se),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(address[1]),
	.D(n88),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[2]  (
	.SI(current_state[1]),
	.SE(test_se),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(current_state[2]),
	.D(n92),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[0]  (
	.SI(n17),
	.SE(test_se),
	.RN(rst_n),
	.Q(current_state[0]),
	.D(n94),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[3]  (
	.SI(current_state[2]),
	.SE(test_se),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(current_state[3]),
	.D(n93),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[1]  (
	.SI(n97),
	.SE(test_se),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(current_state[1]),
	.D(n91),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \address_reg[2]  (
	.SI(address[1]),
	.SE(test_se),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.QN(n18),
	.Q(address[2]),
	.D(n89),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \address_reg[3]  (
	.SI(address[2]),
	.SE(test_se),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.QN(n17),
	.Q(FE_OFN12_address_3_),
	.D(n90),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \address_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(rst_n),
	.QN(n19),
	.Q(address[0]),
	.D(n87),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U16 (
	.Y(alu_fun[2]),
	.B(n23),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U17 (
	.Y(alu_fun[3]),
	.B(n22),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U18 (
	.Y(alu_en),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U19 (
	.Y(n86),
	.B(n46),
	.A(n45), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U20 (
	.Y(n45),
	.B(n96),
	.AN(n60), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U21 (
	.Y(n46),
	.B(n98),
	.AN(n60), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U22 (
	.Y(n60),
	.B(current_state[2]),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U23 (
	.Y(n31),
	.C(n60),
	.B(n100),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U24 (
	.Y(n94),
	.B0(n73),
	.A1(n52),
	.A0(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U25 (
	.Y(n73),
	.B0(n52),
	.A2(n75),
	.A1(n64),
	.A0(n74), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U26 (
	.Y(n74),
	.D(n62),
	.C(n58),
	.B(n81),
	.A(n80), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U27 (
	.Y(n75),
	.B1(n76),
	.B0(n16),
	.A2(n99),
	.A1(n59),
	.A0(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U28 (
	.Y(w_data[0]),
	.B(n25),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U29 (
	.Y(n68),
	.C(n100),
	.B(n97),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U30 (
	.Y(n33),
	.B(n30),
	.AN(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U31 (
	.Y(n93),
	.C0(n20),
	.B0(n62),
	.A1(n16),
	.A0(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U32 (
	.Y(n20),
	.A(n72), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U33 (
	.Y(n72),
	.B0(n99),
	.A2(n50),
	.A1(n52),
	.A0(n59), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U34 (
	.Y(w_data[1]),
	.B(n24),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U35 (
	.Y(w_data[2]),
	.B(n23),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U36 (
	.Y(w_data[3]),
	.B(n22),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U37 (
	.Y(w_data[4]),
	.B(n21),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U38 (
	.Y(r_en),
	.B(n99),
	.A(n47), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U39 (
	.Y(n15),
	.A(n49), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U40 (
	.Y(n96),
	.A(n79), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U41 (
	.Y(n98),
	.A(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U42 (
	.Y(n47),
	.B(n79),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U43 (
	.Y(n80),
	.C(n34),
	.B(n16),
	.A(n79), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U44 (
	.Y(alu_fun[1]),
	.B(n24),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U45 (
	.Y(alu_fun[0]),
	.B(n25),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U46 (
	.Y(clk_en),
	.C0(n85),
	.B0(n33),
	.A1(n58),
	.A0(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U47 (
	.Y(n85),
	.B0(alu_en),
	.A2(current_state[2]),
	.A1(n99),
	.A0(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U48 (
	.Y(w_en),
	.B0(n29),
	.A2(n28),
	.A1(address[1]),
	.A0(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U49 (
	.Y(n27),
	.C(n18),
	.B(n16),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB2XLM U50 (
	.Y(n28),
	.B1(n19),
	.B0(n30),
	.A1N(n31),
	.A0N(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U51 (
	.Y(n57),
	.C(current_state[2]),
	.B(current_state[1]),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U52 (
	.Y(n30),
	.B(current_state[3]),
	.A(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U53 (
	.Y(n97),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U54 (
	.Y(n100),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U55 (
	.Y(n99),
	.A(current_state[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI33X2M U57 (
	.Y(n48),
	.B2(rx_d_valid),
	.B1(current_state[2]),
	.B0(n51),
	.A2(n50),
	.A1(n16),
	.A0(n34), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U58 (
	.Y(n51),
	.C(current_state[0]),
	.B(current_state[3]),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X2M U59 (
	.Y(n32),
	.B0(n29),
	.A1(n33),
	.A0(rx_d_valid), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U60 (
	.Y(n49),
	.B0(n48),
	.A1(n33),
	.A0(rx_d_valid), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U61 (
	.Y(n87),
	.C1(n49),
	.C0(n19),
	.B1(n31),
	.B0(n15),
	.A1(n25),
	.A0(n48), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U62 (
	.Y(n34),
	.B(current_state[3]),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U63 (
	.Y(n89),
	.B1(n23),
	.B0(n48),
	.A1(n18),
	.A0(n49), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U64 (
	.Y(n90),
	.B1(n22),
	.B0(n48),
	.A1(n17),
	.A0(n49), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U65 (
	.Y(n79),
	.B(current_state[1]),
	.A(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U66 (
	.Y(w_data[5]),
	.B(n32),
	.AN(rx_P_data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U67 (
	.Y(w_data[6]),
	.B(n32),
	.AN(rx_P_data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U68 (
	.Y(w_data[7]),
	.B(n32),
	.AN(rx_P_data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U69 (
	.Y(n50),
	.B(current_state[0]),
	.A(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U70 (
	.Y(tx_P_data[0]),
	.B0(n44),
	.A1N(n26),
	.A0N(rd_data[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U71 (
	.Y(n44),
	.B1(n37),
	.B0(alu_out[0]),
	.A1(n36),
	.A0(alu_out[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U72 (
	.Y(tx_P_data[1]),
	.B0(n43),
	.A1N(n26),
	.A0N(rd_data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U73 (
	.Y(n43),
	.B1(n37),
	.B0(alu_out[1]),
	.A1(n36),
	.A0(alu_out[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U74 (
	.Y(tx_P_data[2]),
	.B0(n42),
	.A1N(n26),
	.A0N(rd_data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U75 (
	.Y(n42),
	.B1(n37),
	.B0(alu_out[2]),
	.A1(n36),
	.A0(alu_out[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U76 (
	.Y(tx_P_data[3]),
	.B0(n41),
	.A1N(n26),
	.A0N(rd_data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U77 (
	.Y(n41),
	.B1(n37),
	.B0(alu_out[3]),
	.A1(n36),
	.A0(alu_out[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U78 (
	.Y(tx_P_data[4]),
	.B0(n40),
	.A1N(n26),
	.A0N(rd_data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U79 (
	.Y(n40),
	.B1(n37),
	.B0(alu_out[4]),
	.A1(n36),
	.A0(alu_out[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U80 (
	.Y(tx_P_data[5]),
	.B0(n39),
	.A1N(n26),
	.A0N(rd_data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U81 (
	.Y(n39),
	.B1(n37),
	.B0(alu_out[5]),
	.A1(n36),
	.A0(alu_out[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U82 (
	.Y(tx_P_data[6]),
	.B0(n38),
	.A1N(n26),
	.A0N(rd_data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U83 (
	.Y(n38),
	.B1(n37),
	.B0(alu_out[6]),
	.A1(n36),
	.A0(alu_out[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U84 (
	.Y(tx_P_data[7]),
	.B0(n35),
	.A1N(n26),
	.A0N(rd_data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U85 (
	.Y(n35),
	.B1(n37),
	.B0(alu_out[7]),
	.A1(n36),
	.A0(alu_out[15]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U86 (
	.Y(n54),
	.C0(n63),
	.B0(n62),
	.A1(n96),
	.A0(n61), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U87 (
	.Y(n61),
	.B1(current_state[3]),
	.B0(n59),
	.A1(n34),
	.A0(rx_d_valid), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U88 (
	.Y(n62),
	.D(n82),
	.C(n68),
	.B(rx_P_data[0]),
	.A(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U89 (
	.Y(n82),
	.C(rx_P_data[1]),
	.B(rx_P_data[5]),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U90 (
	.Y(n59),
	.B(full_flag),
	.AN(out_valid), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U91 (
	.Y(n88),
	.B1(n24),
	.B0(n48),
	.A1N(address[1]),
	.A0N(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U92 (
	.Y(n64),
	.B0(n78),
	.A1(n57),
	.A0(rx_d_valid), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B1X2M U93 (
	.Y(n78),
	.B0(n47),
	.A1N(rd_data_valid),
	.A0(full_flag), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U94 (
	.Y(n63),
	.D(n69),
	.C(n68),
	.B(n25),
	.A(n67), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U95 (
	.Y(n69),
	.C(rx_P_data[4]),
	.B(rx_P_data[5]),
	.A(rx_P_data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U96 (
	.Y(n91),
	.B0(n53),
	.A1(n52),
	.A0(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U97 (
	.Y(n53),
	.B0(n52),
	.A2(n56),
	.A1(n55),
	.A0(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U98 (
	.Y(n56),
	.B0(rx_d_valid),
	.A1(n58),
	.A0(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U99 (
	.Y(n55),
	.B0(n98),
	.A1(n60),
	.A0(n59), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U100 (
	.Y(n16),
	.A(rx_d_valid), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U101 (
	.Y(n29),
	.C(n34),
	.B(current_state[1]),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U102 (
	.Y(w_inc),
	.B0(n26),
	.A1(out_valid),
	.A0(alu_en), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U103 (
	.Y(n36),
	.B(out_valid),
	.A(n46), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U104 (
	.Y(n37),
	.B(out_valid),
	.A(n45), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U105 (
	.Y(n26),
	.B(r_en),
	.A(rd_data_valid), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U106 (
	.Y(n58),
	.C(current_state[0]),
	.B(current_state[3]),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U107 (
	.Y(n52),
	.B(current_state[3]),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U108 (
	.Y(n67),
	.C(n83),
	.B(rx_P_data[6]),
	.A(rx_P_data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U109 (
	.Y(n70),
	.C(n83),
	.B(rx_P_data[5]),
	.A(rx_P_data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U110 (
	.Y(n76),
	.B0(n97),
	.A1(n77),
	.A0(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U111 (
	.Y(n77),
	.B(current_state[1]),
	.A(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U112 (
	.Y(n81),
	.D(n84),
	.C(n70),
	.B(n25),
	.A(n68), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U113 (
	.Y(n84),
	.C(rx_P_data[4]),
	.B(rx_P_data[6]),
	.A(rx_P_data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U114 (
	.Y(n25),
	.A(rx_P_data[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U115 (
	.Y(n92),
	.D(n63),
	.C(n66),
	.B(n65),
	.AN(n64), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U116 (
	.Y(n65),
	.B0(current_state[2]),
	.A1N(current_state[0]),
	.A0N(n52), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U117 (
	.Y(n66),
	.D(n71),
	.C(n70),
	.B(rx_P_data[0]),
	.A(n68), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U118 (
	.Y(n71),
	.C(rx_P_data[2]),
	.B(rx_P_data[6]),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U119 (
	.Y(n21),
	.A(rx_P_data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U120 (
	.Y(n24),
	.A(rx_P_data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U121 (
	.Y(n23),
	.A(rx_P_data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U122 (
	.Y(n22),
	.A(rx_P_data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U123 (
	.Y(n83),
	.C(rx_d_valid),
	.B(rx_P_data[3]),
	.A(rx_P_data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(clk_div_en),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module data_sync_top_module_test_1 (
	dest_clk, 
	dest_rst_n, 
	unsync_bus, 
	bus_enable, 
	sync_bus, 
	enable_pulse, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input dest_clk;
   input dest_rst_n;
   input [7:0] unsync_bus;
   input bus_enable;
   output [7:0] sync_bus;
   output enable_pulse;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire sync_bus_enable;
   wire mux_enable;
   wire n1;
   wire n2;

   // Module instantiations
   enable_sync_test_1 dut1 (
	.clk(dest_clk),
	.rst_n(dest_rst_n),
	.bus_enable(bus_enable),
	.sync_bus_enable(sync_bus_enable),
	.test_si(test_si),
	.test_so(n2),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   pulse_gen_test_0 dut2 (
	.clk(dest_clk),
	.rst_n(dest_rst_n),
	.in(sync_bus_enable),
	.d2(mux_enable),
	.out(enable_pulse),
	.test_si(n2),
	.test_so(n1),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   enabled_ff_test_1 dut3 (
	.unsync_bus({ unsync_bus[7],
		unsync_bus[6],
		unsync_bus[5],
		unsync_bus[4],
		unsync_bus[3],
		unsync_bus[2],
		unsync_bus[1],
		unsync_bus[0] }),
	.enable_signal(mux_enable),
	.clk(dest_clk),
	.rst_n(dest_rst_n),
	.sync_bus({ sync_bus[7],
		sync_bus[6],
		sync_bus[5],
		sync_bus[4],
		sync_bus[3],
		sync_bus[2],
		sync_bus[1],
		sync_bus[0] }),
	.test_si(n1),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module enable_sync_test_1 (
	clk, 
	rst_n, 
	bus_enable, 
	sync_bus_enable, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input clk;
   input rst_n;
   input bus_enable;
   output sync_bus_enable;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \enable_sync_reg[1] ;

   assign test_so = \enable_sync_reg[1]  ;

   // Module instantiations
   SDFFRQX2M \enable_sync_reg_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(rst_n),
	.Q(sync_bus_enable),
	.D(\enable_sync_reg[1] ),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \enable_sync_reg_reg[1]  (
	.SI(sync_bus_enable),
	.SE(test_se),
	.RN(rst_n),
	.Q(\enable_sync_reg[1] ),
	.D(bus_enable),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module pulse_gen_test_0 (
	clk, 
	rst_n, 
	in, 
	d2, 
	out, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input clk;
   input rst_n;
   input in;
   output d2;
   output out;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire q;

   assign test_so = q ;

   // Module instantiations
   SDFFRQX2M q_reg (
	.SI(out),
	.SE(test_se),
	.RN(rst_n),
	.Q(q),
	.D(in),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M out_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(rst_n),
	.Q(out),
	.D(d2),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U5 (
	.Y(d2),
	.B(q),
	.AN(in), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module enabled_ff_test_1 (
	unsync_bus, 
	enable_signal, 
	clk, 
	rst_n, 
	sync_bus, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input [7:0] unsync_bus;
   input enable_signal;
   input clk;
   input rst_n;
   output [7:0] sync_bus;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n3;
   wire n5;
   wire n7;
   wire n9;
   wire n11;
   wire n13;
   wire n15;
   wire n17;
   wire n1;

   // Module instantiations
   SDFFRQX2M \sync_bus_reg[7]  (
	.SI(sync_bus[6]),
	.SE(test_se),
	.RN(rst_n),
	.Q(sync_bus[7]),
	.D(n17),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[3]  (
	.SI(sync_bus[2]),
	.SE(test_se),
	.RN(rst_n),
	.Q(sync_bus[3]),
	.D(n9),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[6]  (
	.SI(sync_bus[5]),
	.SE(test_se),
	.RN(rst_n),
	.Q(sync_bus[6]),
	.D(n15),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[5]  (
	.SI(sync_bus[4]),
	.SE(test_se),
	.RN(rst_n),
	.Q(sync_bus[5]),
	.D(n13),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(rst_n),
	.Q(sync_bus[0]),
	.D(n3),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[4]  (
	.SI(sync_bus[3]),
	.SE(test_se),
	.RN(rst_n),
	.Q(sync_bus[4]),
	.D(n11),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[2]  (
	.SI(sync_bus[1]),
	.SE(test_se),
	.RN(rst_n),
	.Q(sync_bus[2]),
	.D(n7),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[1]  (
	.SI(sync_bus[0]),
	.SE(test_se),
	.RN(rst_n),
	.Q(sync_bus[1]),
	.D(n5),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U2 (
	.Y(n1),
	.A(enable_signal), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U3 (
	.Y(n3),
	.B1(n1),
	.B0(sync_bus[0]),
	.A1(enable_signal),
	.A0(unsync_bus[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U4 (
	.Y(n5),
	.B1(n1),
	.B0(sync_bus[1]),
	.A1(enable_signal),
	.A0(unsync_bus[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U5 (
	.Y(n7),
	.B1(n1),
	.B0(sync_bus[2]),
	.A1(enable_signal),
	.A0(unsync_bus[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U6 (
	.Y(n9),
	.B1(n1),
	.B0(sync_bus[3]),
	.A1(enable_signal),
	.A0(unsync_bus[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U7 (
	.Y(n11),
	.B1(n1),
	.B0(sync_bus[4]),
	.A1(enable_signal),
	.A0(unsync_bus[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U8 (
	.Y(n13),
	.B1(n1),
	.B0(sync_bus[5]),
	.A1(enable_signal),
	.A0(unsync_bus[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U9 (
	.Y(n15),
	.B1(n1),
	.B0(sync_bus[6]),
	.A1(enable_signal),
	.A0(unsync_bus[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U10 (
	.Y(n17),
	.B1(n1),
	.B0(sync_bus[7]),
	.A1(enable_signal),
	.A0(unsync_bus[7]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module RX_TOP_MODULE_test_1 (
	rx_in, 
	prescale, 
	parity_enable, 
	parity_type, 
	rx_clk, 
	rst_n, 
	p_data, 
	stop_error, 
	parity_error, 
	start_glitch, 
	data_valid, 
	test_si2, 
	test_si1, 
	test_se, 
	n23, 
	FE_PT1_n24, 
	VDD, 
	VSS);
   input rx_in;
   input [5:0] prescale;
   input parity_enable;
   input parity_type;
   input rx_clk;
   input rst_n;
   output [7:0] p_data;
   output stop_error;
   output parity_error;
   output start_glitch;
   output data_valid;
   input test_si2;
   input test_si1;
   input test_se;
   input n23;
   input FE_PT1_n24;
   inout VDD;
   inout VSS;

   // Internal wires
   wire data_sampler_enable;
   wire sampling_tick;
   wire sampled_bit;
   wire counter_enable;
   wire deserializer_enable;
   wire edge_done_tick;
   wire data_done_tick;
   wire parity_check_enable;
   wire start_check_enable;
   wire stop_check_enable;
   wire n3;
   wire n4;
   wire n5;
   wire n6;

   // Module instantiations
   data_sampler_test_1 dut0 (
	.rx_clk(rx_clk),
	.rst_n(rst_n),
	.data_sampler_enable(data_sampler_enable),
	.sampling_tick(sampling_tick),
	.rx_in(rx_in),
	.sampled_bit(sampled_bit),
	.test_si(test_si1),
	.test_so(n6),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   edge_bit_counter_test_1 dut1 (
	.rx_clk(rx_clk),
	.rst_n(rst_n),
	.prescale({ prescale[5],
		prescale[4],
		prescale[3],
		prescale[2],
		prescale[1],
		prescale[0] }),
	.counter_enable(counter_enable),
	.deserializer_enable(deserializer_enable),
	.edge_done_tick(edge_done_tick),
	.data_done_tick(data_done_tick),
	.sampling_tick(sampling_tick),
	.test_si(n6),
	.test_so(n5),
	.test_se(test_se),
	.n23(n23),
	.FE_PT1_n24(FE_PT1_n24), 
	.VDD(VDD), 
	.VSS(VSS));
   fsm_test_1 dut2 (
	.rx_clk(rx_clk),
	.rst_n(rst_n),
	.rx_in(rx_in),
	.parity_enable(parity_enable),
	.edge_done_tick(edge_done_tick),
	.data_done_tick(data_done_tick),
	.parity_error(parity_error),
	.start_glitch(start_glitch),
	.stop_error(stop_error),
	.deserializer_enable(deserializer_enable),
	.data_sampler_enable(data_sampler_enable),
	.parity_check_enable(parity_check_enable),
	.start_check_enable(start_check_enable),
	.stop_check_enable(stop_check_enable),
	.counter_enable(counter_enable),
	.data_valid(data_valid),
	.test_si(n5),
	.test_so(n4),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   deserializer_test_1 dut3 (
	.sampled_bit(sampled_bit),
	.rx_clk(rx_clk),
	.rst_n(rst_n),
	.deserializer_enable(deserializer_enable),
	.p_data({ p_data[7],
		p_data[6],
		p_data[5],
		p_data[4],
		p_data[3],
		p_data[2],
		p_data[1],
		p_data[0] }),
	.test_si(n4),
	.test_so(n3),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   parity_check_test_1 dut4 (
	.parity_check_enable(parity_check_enable),
	.parity_type(parity_type),
	.rx_clk(rx_clk),
	.rst_n(rst_n),
	.sampled_bit(sampled_bit),
	.p_data({ p_data[7],
		p_data[6],
		p_data[5],
		p_data[4],
		p_data[3],
		p_data[2],
		p_data[1],
		p_data[0] }),
	.parity_error(parity_error),
	.test_si(n3),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   start_check dut5 (
	.start_check_enable(start_check_enable),
	.sampled_bit(sampled_bit),
	.start_glitch(start_glitch), 
	.VDD(VDD), 
	.VSS(VSS));
   stop_check_test_1 dut6 (
	.stop_check_enable(stop_check_enable),
	.rx_clk(rx_clk),
	.rst_n(rst_n),
	.sampled_bit(sampled_bit),
	.stop_error(stop_error),
	.test_si(test_si2),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module data_sampler_test_1 (
	rx_clk, 
	rst_n, 
	data_sampler_enable, 
	sampling_tick, 
	rx_in, 
	sampled_bit, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input rx_clk;
   input rst_n;
   input data_sampler_enable;
   input sampling_tick;
   input rx_in;
   output sampled_bit;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n3;
   wire n7;
   wire n9;
   wire n11;
   wire n13;
   wire n15;
   wire n2;
   wire n4;
   wire n5;
   wire n6;
   wire [2:0] sampled_data;

   assign test_so = n4 ;

   // Module instantiations
   SDFFRQX2M \sampled_data_reg[2]  (
	.SI(n5),
	.SE(test_se),
	.RN(rst_n),
	.Q(sampled_data[2]),
	.D(n15),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sampled_data_reg[0]  (
	.SI(sampled_bit),
	.SE(test_se),
	.RN(rst_n),
	.Q(sampled_data[0]),
	.D(n11),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sampled_data_reg[1]  (
	.SI(sampled_data[0]),
	.SE(test_se),
	.RN(rst_n),
	.Q(sampled_data[1]),
	.D(n13),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M sampled_bit_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(rst_n),
	.Q(sampled_bit),
	.D(n9),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U2 (
	.Y(n11),
	.B1(n5),
	.B0(n7),
	.A1(n6),
	.A0(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U3 (
	.Y(n13),
	.B1(n4),
	.B0(n7),
	.A1(n5),
	.A0(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U4 (
	.Y(n2),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U5 (
	.Y(n7),
	.B(data_sampler_enable),
	.A(sampling_tick), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U6 (
	.Y(n15),
	.B1(n4),
	.B0(n2),
	.A1N(n2),
	.A0N(rx_in), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U7 (
	.Y(n9),
	.B1(n2),
	.B0(n1),
	.A1N(n2),
	.A0N(sampled_bit), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U8 (
	.Y(n1),
	.B0(n3),
	.A1(sampled_data[0]),
	.A0(sampled_data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U9 (
	.Y(n3),
	.B0(n4),
	.A1(n6),
	.A0(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U10 (
	.Y(n5),
	.A(sampled_data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U11 (
	.Y(n4),
	.A(sampled_data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U12 (
	.Y(n6),
	.A(sampled_data[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module edge_bit_counter_test_1 (
	rx_clk, 
	rst_n, 
	prescale, 
	counter_enable, 
	deserializer_enable, 
	edge_done_tick, 
	data_done_tick, 
	sampling_tick, 
	test_si, 
	test_so, 
	test_se, 
	n23, 
	FE_PT1_n24, 
	VDD, 
	VSS);
   input rx_clk;
   input rst_n;
   input [5:0] prescale;
   input counter_enable;
   input deserializer_enable;
   output edge_done_tick;
   output data_done_tick;
   output sampling_tick;
   input test_si;
   output test_so;
   input test_se;
   input n23;
   input FE_PT1_n24;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N4;
   wire N5;
   wire N6;
   wire N7;
   wire N8;
   wire N9;
   wire N12;
   wire N13;
   wire N14;
   wire N15;
   wire N16;
   wire N17;
   wire N19;
   wire N20;
   wire N21;
   wire N22;
   wire N23;
   wire N29;
   wire N30;
   wire N31;
   wire N32;
   wire N33;
   wire N34;
   wire N35;
   wire N36;
   wire N37;
   wire N38;
   wire N39;
   wire N40;
   wire n34;
   wire n35;
   wire n36;
   wire \add_24/carry[5] ;
   wire \add_24/carry[4] ;
   wire \add_24/carry[3] ;
   wire \add_24/carry[2] ;
   wire \add_17/carry[4] ;
   wire \add_17/carry[3] ;
   wire \add_17/carry[2] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire [5:0] edge_counter;
   wire [2:0] data_bit_counter;

   assign test_so = edge_counter[5] ;

   // Module instantiations
   SDFFRQX2M \data_bit_counter_reg[2]  (
	.SI(data_bit_counter[1]),
	.SE(test_se),
	.RN(rst_n),
	.Q(data_bit_counter[2]),
	.D(n35),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \data_bit_counter_reg[1]  (
	.SI(data_bit_counter[0]),
	.SE(test_se),
	.RN(rst_n),
	.Q(data_bit_counter[1]),
	.D(n34),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \data_bit_counter_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(rst_n),
	.Q(data_bit_counter[0]),
	.D(n36),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_counter_reg[5]  (
	.SI(edge_counter[4]),
	.SE(test_se),
	.RN(rst_n),
	.Q(edge_counter[5]),
	.D(N40),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_counter_reg[0]  (
	.SI(data_bit_counter[2]),
	.SE(test_se),
	.RN(rst_n),
	.Q(edge_counter[0]),
	.D(N35),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_counter_reg[4]  (
	.SI(edge_counter[3]),
	.SE(test_se),
	.RN(rst_n),
	.Q(edge_counter[4]),
	.D(N39),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_counter_reg[3]  (
	.SI(edge_counter[2]),
	.SE(test_se),
	.RN(rst_n),
	.Q(edge_counter[3]),
	.D(N38),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_counter_reg[2]  (
	.SI(edge_counter[1]),
	.SE(test_se),
	.RN(rst_n),
	.Q(edge_counter[2]),
	.D(N37),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_counter_reg[1]  (
	.SI(N29),
	.SE(test_se),
	.RN(rst_n),
	.Q(edge_counter[1]),
	.D(N36),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U6 (
	.Y(n1),
	.B(prescale[0]),
	.A(prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U7 (
	.Y(n5),
	.B(prescale[1]),
	.A(prescale[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U8 (
	.S(N21),
	.CO(\add_17/carry[4] ),
	.B(\add_17/carry[3] ),
	.A(prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U9 (
	.S(N20),
	.CO(\add_17/carry[3] ),
	.B(\add_17/carry[2] ),
	.A(prescale[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U10 (
	.S(N19),
	.CO(\add_17/carry[2] ),
	.B(prescale[1]),
	.A(prescale[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U11 (
	.S(N22),
	.CO(N23),
	.B(\add_17/carry[4] ),
	.A(prescale[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U12 (
	.S(N30),
	.CO(\add_24/carry[2] ),
	.B(edge_counter[0]),
	.A(edge_counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U19 (
	.S(N31),
	.CO(\add_24/carry[3] ),
	.B(\add_24/carry[2] ),
	.A(edge_counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U20 (
	.S(N32),
	.CO(\add_24/carry[4] ),
	.B(\add_24/carry[3] ),
	.A(edge_counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U21 (
	.S(N33),
	.CO(\add_24/carry[5] ),
	.B(\add_24/carry[4] ),
	.A(edge_counter[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U23 (
	.Y(N4),
	.B0(n1),
	.A1N(prescale[1]),
	.A0N(prescale[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U24 (
	.Y(n2),
	.B(prescale[2]),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U25 (
	.Y(N5),
	.B0(n2),
	.A1N(prescale[2]),
	.A0N(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U26 (
	.Y(n3),
	.B(prescale[3]),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U27 (
	.Y(N6),
	.B0(n3),
	.A1N(prescale[3]),
	.A0N(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U28 (
	.Y(n4),
	.B(prescale[4]),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U29 (
	.Y(N7),
	.B0(n4),
	.A1N(prescale[4]),
	.A0N(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U30 (
	.Y(N9),
	.B(prescale[5]),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U31 (
	.Y(N8),
	.B0(N9),
	.A1(prescale[5]),
	.A0(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U33 (
	.Y(N12),
	.B0(n5),
	.A1N(prescale[2]),
	.A0N(prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U34 (
	.Y(n6),
	.B(prescale[3]),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U35 (
	.Y(N13),
	.B0(n6),
	.A1N(prescale[3]),
	.A0N(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U36 (
	.Y(N14),
	.B(n6),
	.A(prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X1M U37 (
	.Y(N16),
	.C(n6),
	.B(prescale[5]),
	.A(prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U38 (
	.Y(n7),
	.B0(prescale[5]),
	.A1(n6),
	.A0(prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U39 (
	.Y(N15),
	.B(n7),
	.AN(N16), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U40 (
	.Y(N29),
	.A(edge_counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U41 (
	.Y(N34),
	.B(edge_counter[5]),
	.A(\add_24/carry[5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U42 (
	.Y(n8),
	.B(edge_counter[0]),
	.AN(FE_PT1_n24), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U43 (
	.Y(n12),
	.B1(n8),
	.B0(N4),
	.A1N(edge_counter[1]),
	.A0(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U44 (
	.Y(n11),
	.B(edge_counter[5]),
	.A(N8), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U45 (
	.Y(n9),
	.B(FE_PT1_n24),
	.AN(edge_counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U46 (
	.Y(n10),
	.B1(n9),
	.B0(edge_counter[1]),
	.A1N(N4),
	.A0(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U47 (
	.Y(n25),
	.D(n10),
	.C(n11),
	.B(n12),
	.AN(N9), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U48 (
	.Y(n24),
	.B(edge_counter[4]),
	.A(N7), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U49 (
	.Y(n14),
	.B(edge_counter[2]),
	.A(N5), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U50 (
	.Y(n13),
	.B(edge_counter[3]),
	.A(N6), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U51 (
	.Y(edge_done_tick),
	.D(n13),
	.C(n14),
	.B(n24),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U52 (
	.Y(n26),
	.B(n23),
	.AN(edge_counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U53 (
	.Y(n29),
	.B1(n26),
	.B0(edge_counter[1]),
	.A1N(N12),
	.A0(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U54 (
	.Y(n27),
	.B(edge_counter[0]),
	.AN(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U55 (
	.Y(n28),
	.B1(n27),
	.B0(N12),
	.A1N(edge_counter[1]),
	.A0(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BBX1M U56 (
	.Y(n33),
	.D(n28),
	.C(n29),
	.BN(edge_counter[5]),
	.AN(N16), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U57 (
	.Y(n32),
	.B(edge_counter[4]),
	.A(N15), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U58 (
	.Y(n31),
	.B(edge_counter[2]),
	.A(N13), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U59 (
	.Y(n30),
	.B(edge_counter[3]),
	.A(N14), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U60 (
	.Y(N17),
	.D(n30),
	.C(n31),
	.B(n32),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   OR3X1M U61 (
	.Y(sampling_tick),
	.C(n38),
	.B(n37),
	.A(N17), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U62 (
	.Y(n38),
	.D(n42),
	.C(n41),
	.B(n40),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U63 (
	.Y(n42),
	.B(N23),
	.A(edge_counter[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U64 (
	.Y(n41),
	.B(N21),
	.A(edge_counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U65 (
	.Y(n40),
	.B(N20),
	.A(edge_counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X1M U66 (
	.Y(n39),
	.C(n45),
	.B(n44),
	.A(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U67 (
	.Y(n45),
	.B(n23),
	.A(edge_counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U68 (
	.Y(n44),
	.B(N19),
	.A(edge_counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U69 (
	.Y(n43),
	.B(N22),
	.A(edge_counter[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U70 (
	.Y(n37),
	.D(n48),
	.C(edge_counter[5]),
	.B(n47),
	.A(n46), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U71 (
	.Y(n48),
	.B(edge_counter[0]),
	.A(prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U72 (
	.Y(n47),
	.B(edge_counter[4]),
	.A(prescale[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X1M U73 (
	.Y(n46),
	.C(n51),
	.B(n50),
	.A(n49), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U74 (
	.Y(n51),
	.B(prescale[3]),
	.A(edge_counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U75 (
	.Y(n50),
	.B(prescale[4]),
	.A(edge_counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U76 (
	.Y(n49),
	.B(prescale[2]),
	.A(edge_counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U77 (
	.Y(n36),
	.B(data_bit_counter[0]),
	.A(n52), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U78 (
	.Y(n35),
	.A(n53), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U79 (
	.Y(n53),
	.B1(data_bit_counter[2]),
	.B0(n55),
	.A2(data_bit_counter[1]),
	.A1(data_bit_counter[0]),
	.A0(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U80 (
	.Y(n55),
	.B(n57),
	.A(n56), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U81 (
	.Y(n34),
	.S0(data_bit_counter[1]),
	.B(n57),
	.A(n58), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U82 (
	.Y(n57),
	.B(n52),
	.A(data_bit_counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U83 (
	.Y(n52),
	.B0(n56),
	.A1(n60),
	.A0(n59), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U84 (
	.Y(n58),
	.B(data_bit_counter[0]),
	.A(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U85 (
	.Y(n54),
	.A(n56), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U86 (
	.Y(n56),
	.D(n59),
	.C(edge_done_tick),
	.B(counter_enable),
	.A(deserializer_enable), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U87 (
	.Y(data_done_tick),
	.A(n59), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X1M U88 (
	.Y(n59),
	.C(data_bit_counter[2]),
	.B(data_bit_counter[0]),
	.A(data_bit_counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U89 (
	.Y(N40),
	.B(n61),
	.AN(N34), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U90 (
	.Y(N39),
	.B(n61),
	.AN(N33), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U91 (
	.Y(N38),
	.B(n61),
	.AN(N32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U92 (
	.Y(N37),
	.B(n61),
	.AN(N31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U93 (
	.Y(N36),
	.B(n61),
	.AN(N30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U94 (
	.Y(N35),
	.B(n61),
	.AN(N29), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U95 (
	.Y(n61),
	.B(n60),
	.A(counter_enable), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U96 (
	.Y(n60),
	.A(edge_done_tick), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module fsm_test_1 (
	rx_clk, 
	rst_n, 
	rx_in, 
	parity_enable, 
	edge_done_tick, 
	data_done_tick, 
	parity_error, 
	start_glitch, 
	stop_error, 
	deserializer_enable, 
	data_sampler_enable, 
	parity_check_enable, 
	start_check_enable, 
	stop_check_enable, 
	counter_enable, 
	data_valid, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input rx_clk;
   input rst_n;
   input rx_in;
   input parity_enable;
   input edge_done_tick;
   input data_done_tick;
   input parity_error;
   input start_glitch;
   input stop_error;
   output deserializer_enable;
   output data_sampler_enable;
   output parity_check_enable;
   output start_check_enable;
   output stop_check_enable;
   output counter_enable;
   output data_valid;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire [2:0] current_state;
   wire [2:0] next_state;

   assign test_so = n7 ;

   // Module instantiations
   SDFFRQX2M \current_state_reg[2]  (
	.SI(n9),
	.SE(test_se),
	.RN(rst_n),
	.Q(current_state[2]),
	.D(next_state[2]),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[1]  (
	.SI(current_state[0]),
	.SE(test_se),
	.RN(rst_n),
	.Q(current_state[1]),
	.D(next_state[1]),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(rst_n),
	.Q(current_state[0]),
	.D(next_state[0]),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4XLM U6 (
	.Y(data_valid),
	.D(n15),
	.C(n5),
	.B(parity_error),
	.A(stop_error), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U7 (
	.Y(n13),
	.B(n7),
	.A(edge_done_tick), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U8 (
	.Y(n21),
	.B0(n14),
	.A1(n5),
	.A0(start_glitch), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U9 (
	.Y(n10),
	.A(edge_done_tick), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U10 (
	.Y(parity_check_enable),
	.B(n14),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U11 (
	.Y(next_state[1]),
	.B1(n4),
	.B0(start_glitch),
	.A2(n17),
	.A1(current_state[2]),
	.A0(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U12 (
	.Y(n17),
	.B(n10),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U13 (
	.Y(n4),
	.A(start_check_enable), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U14 (
	.Y(n18),
	.B0(current_state[0]),
	.A1(n11),
	.A0(data_done_tick), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U15 (
	.Y(deserializer_enable),
	.C(n9),
	.B(current_state[0]),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U16 (
	.Y(start_check_enable),
	.C(n5),
	.B(current_state[1]),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U17 (
	.Y(next_state[0]),
	.C0(n20),
	.B0(n19),
	.A1(counter_enable),
	.A0(rx_in), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U18 (
	.Y(n19),
	.C(parity_enable),
	.B(data_done_tick),
	.A(deserializer_enable), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI33XLM U19 (
	.Y(n20),
	.B2(n21),
	.B1(n10),
	.B0(n7),
	.A2(n8),
	.A1(n5),
	.A0(edge_done_tick), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n8),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U21 (
	.Y(next_state[2]),
	.B1(n13),
	.B0(n16),
	.A1(n15),
	.A0(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U22 (
	.Y(n16),
	.B0(n6),
	.A2(data_done_tick),
	.A1(n11),
	.A0(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U23 (
	.Y(n6),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3BX2M U24 (
	.Y(stop_check_enable),
	.C(n7),
	.B(n10),
	.AN(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U25 (
	.Y(n5),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U26 (
	.Y(data_sampler_enable),
	.B(n7),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U27 (
	.Y(n9),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U28 (
	.Y(n7),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U29 (
	.Y(counter_enable),
	.B(n9),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U30 (
	.Y(n22),
	.B(current_state[0]),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U31 (
	.Y(n14),
	.B(current_state[0]),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U32 (
	.Y(n15),
	.B(n9),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U33 (
	.Y(n12),
	.B(current_state[1]),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U34 (
	.Y(n11),
	.A(parity_enable), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module deserializer_test_1 (
	sampled_bit, 
	rx_clk, 
	rst_n, 
	deserializer_enable, 
	p_data, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input sampled_bit;
   input rx_clk;
   input rst_n;
   input deserializer_enable;
   output [7:0] p_data;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n10;
   wire n12;
   wire n14;
   wire n16;
   wire n18;
   wire n20;
   wire n22;
   wire n24;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n25;

   assign test_so = n2 ;

   // Module instantiations
   SDFFRQX2M \p_data_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(rst_n),
	.Q(p_data[0]),
	.D(n10),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \p_data_reg[7]  (
	.SI(n3),
	.SE(test_se),
	.RN(rst_n),
	.Q(p_data[7]),
	.D(n24),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \p_data_reg[3]  (
	.SI(n7),
	.SE(test_se),
	.RN(rst_n),
	.Q(p_data[3]),
	.D(n16),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \p_data_reg[6]  (
	.SI(n4),
	.SE(test_se),
	.RN(rst_n),
	.Q(p_data[6]),
	.D(n22),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \p_data_reg[5]  (
	.SI(n5),
	.SE(test_se),
	.RN(rst_n),
	.Q(p_data[5]),
	.D(n20),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \p_data_reg[2]  (
	.SI(n8),
	.SE(test_se),
	.RN(rst_n),
	.Q(p_data[2]),
	.D(n14),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \p_data_reg[4]  (
	.SI(n6),
	.SE(test_se),
	.RN(rst_n),
	.Q(p_data[4]),
	.D(n18),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \p_data_reg[1]  (
	.SI(p_data[0]),
	.SE(test_se),
	.RN(rst_n),
	.Q(p_data[1]),
	.D(n12),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U2 (
	.Y(n25),
	.A(deserializer_enable), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U4 (
	.Y(n12),
	.B1(n8),
	.B0(deserializer_enable),
	.A1(n7),
	.A0(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U5 (
	.Y(n14),
	.B1(n7),
	.B0(deserializer_enable),
	.A1(n6),
	.A0(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U6 (
	.Y(n16),
	.B1(n6),
	.B0(deserializer_enable),
	.A1(n5),
	.A0(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U7 (
	.Y(n18),
	.B1(n5),
	.B0(deserializer_enable),
	.A1(n4),
	.A0(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U8 (
	.Y(n20),
	.B1(n4),
	.B0(deserializer_enable),
	.A1(n3),
	.A0(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U9 (
	.Y(n22),
	.B1(n3),
	.B0(deserializer_enable),
	.A1(n2),
	.A0(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U10 (
	.Y(n10),
	.B1(n8),
	.B0(n25),
	.A1N(n25),
	.A0N(p_data[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U11 (
	.Y(n24),
	.B1(n2),
	.B0(deserializer_enable),
	.A1N(deserializer_enable),
	.A0N(sampled_bit), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U12 (
	.Y(n8),
	.A(p_data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U13 (
	.Y(n5),
	.A(p_data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U14 (
	.Y(n7),
	.A(p_data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U15 (
	.Y(n4),
	.A(p_data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U16 (
	.Y(n3),
	.A(p_data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U17 (
	.Y(n6),
	.A(p_data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U26 (
	.Y(n2),
	.A(p_data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module parity_check_test_1 (
	parity_check_enable, 
	parity_type, 
	rx_clk, 
	rst_n, 
	sampled_bit, 
	p_data, 
	parity_error, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input parity_check_enable;
   input parity_type;
   input rx_clk;
   input rst_n;
   input sampled_bit;
   input [7:0] p_data;
   output parity_error;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n11;
   wire n1;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n9;
   wire n10;
   wire n2;

   // Module instantiations
   OAI2BB2X1M U4 (
	.Y(n9),
	.B1(n10),
	.B0(n1),
	.A1N(n10),
	.A0N(parity_error), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U5 (
	.Y(n1),
	.C(n5),
	.B(n4),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U6 (
	.Y(n10),
	.A(parity_check_enable), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U7 (
	.Y(n5),
	.B(p_data[1]),
	.A(p_data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U8 (
	.Y(n4),
	.C(n6),
	.B(p_data[6]),
	.A(p_data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U9 (
	.Y(n6),
	.B(parity_type),
	.A(sampled_bit), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U10 (
	.Y(n3),
	.C(n7),
	.B(p_data[0]),
	.A(p_data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U12 (
	.Y(n7),
	.B(p_data[4]),
	.A(p_data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M parity_error_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(rst_n),
	.Q(n11),
	.D(n9),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U3 (
	.Y(n2),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX12M U11 (
	.Y(parity_error),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module start_check (
	start_check_enable, 
	sampled_bit, 
	start_glitch, 
	VDD, 
	VSS);
   input start_check_enable;
   input sampled_bit;
   output start_glitch;
   inout VDD;
   inout VSS;

   // Module instantiations
   AND2X12M U3 (
	.Y(start_glitch),
	.B(sampled_bit),
	.A(start_check_enable), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module stop_check_test_1 (
	stop_check_enable, 
	rx_clk, 
	rst_n, 
	sampled_bit, 
	stop_error, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input stop_check_enable;
   input rx_clk;
   input rst_n;
   input sampled_bit;
   output stop_error;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n5;
   wire n3;
   wire n4;
   wire n7;
   wire n8;
   wire n1;

   // Module instantiations
   OAI2BB2X1M U4 (
	.Y(n3),
	.B1(n4),
	.B0(sampled_bit),
	.A1N(n4),
	.A0N(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U6 (
	.Y(n4),
	.A(stop_check_enable), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U8 (
	.Y(n8),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M stop_error_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(rst_n),
	.QN(n7),
	.Q(n5),
	.D(n3),
	.CK(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U3 (
	.Y(n1),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX12M U5 (
	.Y(stop_error),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module RF_test_1 (
	wren, 
	rden, 
	clk, 
	rst, 
	wrdata, 
	address, 
	rddata, 
	rddata_valid, 
	reg0, 
	reg1, 
	reg2, 
	reg3, 
	test_si3, 
	test_si2, 
	test_si1, 
	test_so2, 
	test_so1, 
	test_se, 
	FE_OFN0_scan_rst_sync1_mux_out, 
	FE_OFN2_scan_rst_sync1_mux_out, 
	scan_clk_ref_clk_mux_out__L4_N1, 
	VDD, 
	VSS);
   input wren;
   input rden;
   input clk;
   input rst;
   input [7:0] wrdata;
   input [3:0] address;
   output [7:0] rddata;
   output rddata_valid;
   output [7:0] reg0;
   output [7:0] reg1;
   output [7:0] reg2;
   output [7:0] reg3;
   input test_si3;
   input test_si2;
   input test_si1;
   output test_so2;
   output test_so1;
   input test_se;
   input FE_OFN0_scan_rst_sync1_mux_out;
   input FE_OFN2_scan_rst_sync1_mux_out;
   input scan_clk_ref_clk_mux_out__L4_N1;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_OFN19_reg0_7_;
   wire FE_OFN18_reg0_6_;
   wire FE_OFN17_reg0_5_;
   wire FE_OFN16_reg0_4_;
   wire FE_OFN15_reg0_3_;
   wire FE_OFN14_reg1_7_;
   wire FE_OFN11_SO_2_;
   wire FE_OFN10_SO_1_;
   wire FE_OFN5_scan_rst_sync1_mux_out;
   wire FE_OFN1_scan_rst_sync1_mux_out;
   wire N10;
   wire N11;
   wire N12;
   wire N13;
   wire \reg_file[4][7] ;
   wire \reg_file[4][6] ;
   wire \reg_file[4][5] ;
   wire \reg_file[4][4] ;
   wire \reg_file[4][3] ;
   wire \reg_file[4][2] ;
   wire \reg_file[4][1] ;
   wire \reg_file[4][0] ;
   wire \reg_file[5][7] ;
   wire \reg_file[5][6] ;
   wire \reg_file[5][5] ;
   wire \reg_file[5][4] ;
   wire \reg_file[5][3] ;
   wire \reg_file[5][2] ;
   wire \reg_file[5][1] ;
   wire \reg_file[5][0] ;
   wire \reg_file[6][7] ;
   wire \reg_file[6][6] ;
   wire \reg_file[6][5] ;
   wire \reg_file[6][4] ;
   wire \reg_file[6][3] ;
   wire \reg_file[6][2] ;
   wire \reg_file[6][1] ;
   wire \reg_file[6][0] ;
   wire \reg_file[7][7] ;
   wire \reg_file[7][6] ;
   wire \reg_file[7][5] ;
   wire \reg_file[7][4] ;
   wire \reg_file[7][3] ;
   wire \reg_file[7][2] ;
   wire \reg_file[7][1] ;
   wire \reg_file[7][0] ;
   wire \reg_file[8][7] ;
   wire \reg_file[8][6] ;
   wire \reg_file[8][5] ;
   wire \reg_file[8][4] ;
   wire \reg_file[8][3] ;
   wire \reg_file[8][2] ;
   wire \reg_file[8][1] ;
   wire \reg_file[8][0] ;
   wire \reg_file[9][7] ;
   wire \reg_file[9][6] ;
   wire \reg_file[9][5] ;
   wire \reg_file[9][4] ;
   wire \reg_file[9][3] ;
   wire \reg_file[9][2] ;
   wire \reg_file[9][1] ;
   wire \reg_file[9][0] ;
   wire \reg_file[10][7] ;
   wire \reg_file[10][6] ;
   wire \reg_file[10][5] ;
   wire \reg_file[10][4] ;
   wire \reg_file[10][3] ;
   wire \reg_file[10][2] ;
   wire \reg_file[10][1] ;
   wire \reg_file[10][0] ;
   wire \reg_file[11][7] ;
   wire \reg_file[11][6] ;
   wire \reg_file[11][5] ;
   wire \reg_file[11][4] ;
   wire \reg_file[11][3] ;
   wire \reg_file[11][2] ;
   wire \reg_file[11][1] ;
   wire \reg_file[11][0] ;
   wire \reg_file[12][7] ;
   wire \reg_file[12][6] ;
   wire \reg_file[12][5] ;
   wire \reg_file[12][4] ;
   wire \reg_file[12][3] ;
   wire \reg_file[12][2] ;
   wire \reg_file[12][1] ;
   wire \reg_file[12][0] ;
   wire \reg_file[13][7] ;
   wire \reg_file[13][6] ;
   wire \reg_file[13][5] ;
   wire \reg_file[13][4] ;
   wire \reg_file[13][3] ;
   wire \reg_file[13][2] ;
   wire \reg_file[13][1] ;
   wire \reg_file[13][0] ;
   wire \reg_file[14][7] ;
   wire \reg_file[14][6] ;
   wire \reg_file[14][5] ;
   wire \reg_file[14][4] ;
   wire \reg_file[14][3] ;
   wire \reg_file[14][2] ;
   wire \reg_file[14][1] ;
   wire \reg_file[14][0] ;
   wire \reg_file[15][7] ;
   wire \reg_file[15][6] ;
   wire \reg_file[15][5] ;
   wire \reg_file[15][4] ;
   wire \reg_file[15][3] ;
   wire \reg_file[15][2] ;
   wire \reg_file[15][1] ;
   wire \reg_file[15][0] ;
   wire N35;
   wire N36;
   wire N37;
   wire N38;
   wire N39;
   wire N40;
   wire N41;
   wire N42;
   wire n1;
   wire n2;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n25;
   wire n30;
   wire n31;
   wire n38;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n335;
   wire n336;
   wire n345;
   wire n346;
   wire n347;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;

   assign N10 = address[0] ;
   assign N11 = address[1] ;
   assign N12 = address[2] ;
   assign N13 = address[3] ;
   assign test_so1 = \reg_file[12][5]  ;
   assign test_so2 = \reg_file[15][7]  ;

   // Module instantiations
   BUFX8M FE_OFC19_reg0_7_ (
	.Y(reg0[7]),
	.A(FE_OFN19_reg0_7_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX10M FE_OFC18_reg0_6_ (
	.Y(reg0[6]),
	.A(FE_OFN18_reg0_6_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX10M FE_OFC17_reg0_5_ (
	.Y(reg0[5]),
	.A(FE_OFN17_reg0_5_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX10M FE_OFC16_reg0_4_ (
	.Y(reg0[4]),
	.A(FE_OFN16_reg0_4_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX10M FE_OFC15_reg0_3_ (
	.Y(reg0[3]),
	.A(FE_OFN15_reg0_3_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX8M FE_OFC14_reg1_7_ (
	.Y(reg1[7]),
	.A(FE_OFN14_reg1_7_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX10M FE_OFC11_SO_2_ (
	.Y(reg2[3]),
	.A(FE_OFN11_SO_2_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX10M FE_OFC10_SO_1_ (
	.Y(\reg_file[12][5] ),
	.A(FE_OFN10_SO_1_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX4M FE_OFC5_scan_rst_sync1_mux_out (
	.Y(FE_OFN5_scan_rst_sync1_mux_out),
	.A(FE_OFN1_scan_rst_sync1_mux_out), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX6M FE_OFC1_scan_rst_sync1_mux_out (
	.Y(FE_OFN1_scan_rst_sync1_mux_out),
	.A(FE_OFN0_scan_rst_sync1_mux_out), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \rddata_reg[7]  (
	.SI(rddata[6]),
	.SE(n379),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(rddata[7]),
	.D(n312),
	.CK(scan_clk_ref_clk_mux_out__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \rddata_reg[6]  (
	.SI(rddata[5]),
	.SE(n378),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(rddata[6]),
	.D(n311),
	.CK(scan_clk_ref_clk_mux_out__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \rddata_reg[5]  (
	.SI(rddata[4]),
	.SE(n377),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(rddata[5]),
	.D(n310),
	.CK(scan_clk_ref_clk_mux_out__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \rddata_reg[4]  (
	.SI(rddata[3]),
	.SE(n380),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(rddata[4]),
	.D(n309),
	.CK(scan_clk_ref_clk_mux_out__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \rddata_reg[3]  (
	.SI(rddata[2]),
	.SE(n379),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(rddata[3]),
	.D(n308),
	.CK(scan_clk_ref_clk_mux_out__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \rddata_reg[2]  (
	.SI(rddata[1]),
	.SE(n378),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(rddata[2]),
	.D(n307),
	.CK(scan_clk_ref_clk_mux_out__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \rddata_reg[1]  (
	.SI(rddata[0]),
	.SE(n377),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(rddata[1]),
	.D(n306),
	.CK(scan_clk_ref_clk_mux_out__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \rddata_reg[0]  (
	.SI(test_si1),
	.SE(n380),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(rddata[0]),
	.D(n305),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[5][7]  (
	.SI(\reg_file[5][6] ),
	.SE(n379),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[5][7] ),
	.D(n264),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[5][6]  (
	.SI(\reg_file[5][5] ),
	.SE(n378),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[5][6] ),
	.D(n263),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[5][5]  (
	.SI(\reg_file[5][4] ),
	.SE(n377),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[5][5] ),
	.D(n262),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[5][4]  (
	.SI(\reg_file[5][3] ),
	.SE(n380),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[5][4] ),
	.D(n261),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[5][3]  (
	.SI(\reg_file[5][2] ),
	.SE(n379),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[5][3] ),
	.D(n260),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[5][2]  (
	.SI(\reg_file[5][1] ),
	.SE(n378),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[5][2] ),
	.D(n259),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[5][1]  (
	.SI(\reg_file[5][0] ),
	.SE(n377),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[5][1] ),
	.D(n258),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[5][0]  (
	.SI(\reg_file[4][7] ),
	.SE(n380),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[5][0] ),
	.D(n257),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[9][7]  (
	.SI(\reg_file[9][6] ),
	.SE(n379),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[9][7] ),
	.D(n232),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[9][6]  (
	.SI(\reg_file[9][5] ),
	.SE(n378),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[9][6] ),
	.D(n231),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[9][5]  (
	.SI(\reg_file[9][4] ),
	.SE(n377),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(\reg_file[9][5] ),
	.D(n230),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[9][4]  (
	.SI(\reg_file[9][3] ),
	.SE(n380),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(\reg_file[9][4] ),
	.D(n229),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[9][3]  (
	.SI(\reg_file[9][2] ),
	.SE(n379),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(\reg_file[9][3] ),
	.D(n228),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[9][2]  (
	.SI(\reg_file[9][1] ),
	.SE(n378),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(\reg_file[9][2] ),
	.D(n227),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[9][1]  (
	.SI(\reg_file[9][0] ),
	.SE(n377),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(\reg_file[9][1] ),
	.D(n226),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[9][0]  (
	.SI(\reg_file[8][7] ),
	.SE(n380),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[9][0] ),
	.D(n225),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[13][7]  (
	.SI(\reg_file[13][6] ),
	.SE(n379),
	.RN(rst),
	.Q(\reg_file[13][7] ),
	.D(n200),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[13][6]  (
	.SI(\reg_file[13][5] ),
	.SE(n378),
	.RN(rst),
	.Q(\reg_file[13][6] ),
	.D(n199),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[13][5]  (
	.SI(\reg_file[13][4] ),
	.SE(n377),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(\reg_file[13][5] ),
	.D(n198),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[13][4]  (
	.SI(\reg_file[13][3] ),
	.SE(n380),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(\reg_file[13][4] ),
	.D(n197),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[13][3]  (
	.SI(\reg_file[13][2] ),
	.SE(n379),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(\reg_file[13][3] ),
	.D(n196),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[13][2]  (
	.SI(\reg_file[13][1] ),
	.SE(n378),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(\reg_file[13][2] ),
	.D(n195),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[13][1]  (
	.SI(\reg_file[13][0] ),
	.SE(n377),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(\reg_file[13][1] ),
	.D(n194),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[13][0]  (
	.SI(\reg_file[12][7] ),
	.SE(n380),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(\reg_file[13][0] ),
	.D(n193),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[7][7]  (
	.SI(\reg_file[7][6] ),
	.SE(n379),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[7][7] ),
	.D(n248),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[7][6]  (
	.SI(\reg_file[7][5] ),
	.SE(n378),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[7][6] ),
	.D(n247),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[7][5]  (
	.SI(\reg_file[7][4] ),
	.SE(n377),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[7][5] ),
	.D(n246),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[7][4]  (
	.SI(\reg_file[7][3] ),
	.SE(n380),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[7][4] ),
	.D(n245),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[7][3]  (
	.SI(\reg_file[7][2] ),
	.SE(n379),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[7][3] ),
	.D(n244),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[7][2]  (
	.SI(\reg_file[7][1] ),
	.SE(n378),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[7][2] ),
	.D(n243),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[7][1]  (
	.SI(\reg_file[7][0] ),
	.SE(n377),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[7][1] ),
	.D(n242),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[7][0]  (
	.SI(\reg_file[6][7] ),
	.SE(n380),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[7][0] ),
	.D(n241),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[11][7]  (
	.SI(\reg_file[11][6] ),
	.SE(n379),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[11][7] ),
	.D(n216),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[11][6]  (
	.SI(\reg_file[11][5] ),
	.SE(n378),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[11][6] ),
	.D(n215),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[11][5]  (
	.SI(\reg_file[11][4] ),
	.SE(n377),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[11][5] ),
	.D(n214),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[11][4]  (
	.SI(\reg_file[11][3] ),
	.SE(n380),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[11][4] ),
	.D(n213),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[11][3]  (
	.SI(\reg_file[11][2] ),
	.SE(n379),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(\reg_file[11][3] ),
	.D(n212),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[11][2]  (
	.SI(\reg_file[11][1] ),
	.SE(n378),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(\reg_file[11][2] ),
	.D(n211),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[11][1]  (
	.SI(\reg_file[11][0] ),
	.SE(n377),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(\reg_file[11][1] ),
	.D(n210),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[11][0]  (
	.SI(\reg_file[10][7] ),
	.SE(n380),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(\reg_file[11][0] ),
	.D(n209),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[15][7]  (
	.SI(\reg_file[15][6] ),
	.SE(n379),
	.RN(rst),
	.Q(\reg_file[15][7] ),
	.D(n184),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[15][6]  (
	.SI(\reg_file[15][5] ),
	.SE(n378),
	.RN(rst),
	.Q(\reg_file[15][6] ),
	.D(n183),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[15][5]  (
	.SI(\reg_file[15][4] ),
	.SE(n377),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(\reg_file[15][5] ),
	.D(n182),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[15][4]  (
	.SI(\reg_file[15][3] ),
	.SE(n380),
	.RN(rst),
	.Q(\reg_file[15][4] ),
	.D(n181),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[15][3]  (
	.SI(\reg_file[15][2] ),
	.SE(n379),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(\reg_file[15][3] ),
	.D(n180),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[15][2]  (
	.SI(\reg_file[15][1] ),
	.SE(n378),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(\reg_file[15][2] ),
	.D(n179),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[15][1]  (
	.SI(\reg_file[15][0] ),
	.SE(n377),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(\reg_file[15][1] ),
	.D(n178),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[15][0]  (
	.SI(\reg_file[14][7] ),
	.SE(n380),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[15][0] ),
	.D(n177),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[6][7]  (
	.SI(\reg_file[6][6] ),
	.SE(n379),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[6][7] ),
	.D(n256),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[6][6]  (
	.SI(\reg_file[6][5] ),
	.SE(n378),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[6][6] ),
	.D(n255),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[6][5]  (
	.SI(\reg_file[6][4] ),
	.SE(n377),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[6][5] ),
	.D(n254),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[6][4]  (
	.SI(\reg_file[6][3] ),
	.SE(n380),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[6][4] ),
	.D(n253),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[6][3]  (
	.SI(\reg_file[6][2] ),
	.SE(n379),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[6][3] ),
	.D(n252),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[6][2]  (
	.SI(\reg_file[6][1] ),
	.SE(n378),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[6][2] ),
	.D(n251),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[6][1]  (
	.SI(\reg_file[6][0] ),
	.SE(n377),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[6][1] ),
	.D(n250),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[6][0]  (
	.SI(\reg_file[5][7] ),
	.SE(n380),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[6][0] ),
	.D(n249),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[10][7]  (
	.SI(\reg_file[10][6] ),
	.SE(n379),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[10][7] ),
	.D(n224),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[10][6]  (
	.SI(\reg_file[10][5] ),
	.SE(n378),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[10][6] ),
	.D(n223),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[10][5]  (
	.SI(\reg_file[10][4] ),
	.SE(n377),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[10][5] ),
	.D(n222),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[10][4]  (
	.SI(\reg_file[10][3] ),
	.SE(n380),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(\reg_file[10][4] ),
	.D(n221),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[10][3]  (
	.SI(\reg_file[10][2] ),
	.SE(n379),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(\reg_file[10][3] ),
	.D(n220),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[10][2]  (
	.SI(\reg_file[10][1] ),
	.SE(n378),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(\reg_file[10][2] ),
	.D(n219),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[10][1]  (
	.SI(\reg_file[10][0] ),
	.SE(n377),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(\reg_file[10][1] ),
	.D(n218),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[10][0]  (
	.SI(\reg_file[9][7] ),
	.SE(n380),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[10][0] ),
	.D(n217),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[14][7]  (
	.SI(\reg_file[14][6] ),
	.SE(n379),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[14][7] ),
	.D(n192),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[14][6]  (
	.SI(\reg_file[14][5] ),
	.SE(n378),
	.RN(rst),
	.Q(\reg_file[14][6] ),
	.D(n191),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[14][5]  (
	.SI(\reg_file[14][4] ),
	.SE(n377),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(\reg_file[14][5] ),
	.D(n190),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[14][4]  (
	.SI(\reg_file[14][3] ),
	.SE(n380),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(\reg_file[14][4] ),
	.D(n189),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[14][3]  (
	.SI(\reg_file[14][2] ),
	.SE(n379),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(\reg_file[14][3] ),
	.D(n188),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[14][2]  (
	.SI(\reg_file[14][1] ),
	.SE(n378),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(\reg_file[14][2] ),
	.D(n187),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[14][1]  (
	.SI(\reg_file[14][0] ),
	.SE(n377),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(\reg_file[14][1] ),
	.D(n186),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[14][0]  (
	.SI(\reg_file[13][7] ),
	.SE(n380),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[14][0] ),
	.D(n185),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[4][7]  (
	.SI(\reg_file[4][6] ),
	.SE(n379),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[4][7] ),
	.D(n272),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[4][6]  (
	.SI(\reg_file[4][5] ),
	.SE(n378),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[4][6] ),
	.D(n271),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[4][5]  (
	.SI(\reg_file[4][4] ),
	.SE(n377),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[4][5] ),
	.D(n270),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[4][4]  (
	.SI(\reg_file[4][3] ),
	.SE(n380),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[4][4] ),
	.D(n269),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[4][3]  (
	.SI(\reg_file[4][2] ),
	.SE(n379),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[4][3] ),
	.D(n268),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[4][2]  (
	.SI(\reg_file[4][1] ),
	.SE(n378),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[4][2] ),
	.D(n267),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[4][1]  (
	.SI(\reg_file[4][0] ),
	.SE(n377),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[4][1] ),
	.D(n266),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[4][0]  (
	.SI(reg3[7]),
	.SE(n380),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[4][0] ),
	.D(n265),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[8][7]  (
	.SI(\reg_file[8][6] ),
	.SE(n379),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[8][7] ),
	.D(n240),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[8][6]  (
	.SI(\reg_file[8][5] ),
	.SE(n378),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[8][6] ),
	.D(n239),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[8][5]  (
	.SI(\reg_file[8][4] ),
	.SE(n377),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[8][5] ),
	.D(n238),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[8][4]  (
	.SI(\reg_file[8][3] ),
	.SE(n380),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(\reg_file[8][4] ),
	.D(n237),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[8][3]  (
	.SI(\reg_file[8][2] ),
	.SE(n379),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(\reg_file[8][3] ),
	.D(n236),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[8][2]  (
	.SI(\reg_file[8][1] ),
	.SE(n378),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(\reg_file[8][2] ),
	.D(n235),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[8][1]  (
	.SI(\reg_file[8][0] ),
	.SE(n377),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(\reg_file[8][1] ),
	.D(n234),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[8][0]  (
	.SI(\reg_file[7][7] ),
	.SE(n380),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(\reg_file[8][0] ),
	.D(n233),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[12][7]  (
	.SI(\reg_file[12][6] ),
	.SE(n379),
	.RN(rst),
	.Q(\reg_file[12][7] ),
	.D(n208),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[12][6]  (
	.SI(test_si3),
	.SE(n378),
	.RN(rst),
	.Q(\reg_file[12][6] ),
	.D(n207),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[12][4]  (
	.SI(\reg_file[12][3] ),
	.SE(n380),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(\reg_file[12][4] ),
	.D(n205),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[12][3]  (
	.SI(\reg_file[12][2] ),
	.SE(n379),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(\reg_file[12][3] ),
	.D(n204),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[12][2]  (
	.SI(\reg_file[12][1] ),
	.SE(n378),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(\reg_file[12][2] ),
	.D(n203),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[12][1]  (
	.SI(\reg_file[12][0] ),
	.SE(n377),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(\reg_file[12][1] ),
	.D(n202),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[12][0]  (
	.SI(\reg_file[11][7] ),
	.SE(n380),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(\reg_file[12][0] ),
	.D(n201),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M rddata_valid_reg (
	.SI(rddata[7]),
	.SE(n379),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(rddata_valid),
	.D(n176),
	.CK(scan_clk_ref_clk_mux_out__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX4M \reg_file_reg[1][6]  (
	.SI(reg1[5]),
	.SE(n378),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(reg1[6]),
	.D(n295),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX4M \reg_file_reg[1][1]  (
	.SI(reg1[0]),
	.SE(n377),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(reg1[1]),
	.D(n290),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX2M \reg_file_reg[0][7]  (
	.SI(reg0[6]),
	.SE(n380),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(FE_OFN19_reg0_7_),
	.D(n304),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX4M \reg_file_reg[0][6]  (
	.SI(reg0[5]),
	.SE(n379),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(FE_OFN18_reg0_6_),
	.D(n303),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX2M \reg_file_reg[0][5]  (
	.SI(reg0[4]),
	.SE(n378),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(FE_OFN17_reg0_5_),
	.D(n302),
	.CK(scan_clk_ref_clk_mux_out__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX2M \reg_file_reg[0][4]  (
	.SI(reg0[3]),
	.SE(n377),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(FE_OFN16_reg0_4_),
	.D(n301),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX2M \reg_file_reg[0][3]  (
	.SI(reg0[2]),
	.SE(n380),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(FE_OFN15_reg0_3_),
	.D(n300),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[0][2]  (
	.SI(reg0[1]),
	.SE(n379),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(reg0[2]),
	.D(n299),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[0][1]  (
	.SI(reg0[0]),
	.SE(n378),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(reg0[1]),
	.D(n298),
	.CK(scan_clk_ref_clk_mux_out__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[0][0]  (
	.SI(rddata_valid),
	.SE(n377),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(reg0[0]),
	.D(n297),
	.CK(scan_clk_ref_clk_mux_out__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[2][1]  (
	.SI(reg2[0]),
	.SE(n380),
	.RN(rst),
	.Q(reg2[1]),
	.D(n282),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \reg_file_reg[2][0]  (
	.SN(FE_OFN2_scan_rst_sync1_mux_out),
	.SI(reg1[7]),
	.SE(test_se),
	.Q(reg2[0]),
	.D(n281),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX2M \reg_file_reg[1][7]  (
	.SI(reg1[6]),
	.SE(n379),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(FE_OFN14_reg1_7_),
	.D(n296),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX4M \reg_file_reg[1][5]  (
	.SI(reg1[4]),
	.SE(n378),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(reg1[5]),
	.D(n294),
	.CK(scan_clk_ref_clk_mux_out__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX4M \reg_file_reg[1][4]  (
	.SI(reg1[3]),
	.SE(n377),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(reg1[4]),
	.D(n293),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX4M \reg_file_reg[1][3]  (
	.SI(reg1[2]),
	.SE(n380),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(reg1[3]),
	.D(n292),
	.CK(scan_clk_ref_clk_mux_out__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX4M \reg_file_reg[1][2]  (
	.SI(reg1[1]),
	.SE(n379),
	.RN(FE_OFN5_scan_rst_sync1_mux_out),
	.Q(reg1[2]),
	.D(n291),
	.CK(scan_clk_ref_clk_mux_out__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX4M \reg_file_reg[1][0]  (
	.SI(reg0[7]),
	.SE(n378),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(reg1[0]),
	.D(n289),
	.CK(scan_clk_ref_clk_mux_out__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \reg_file_reg[3][5]  (
	.SN(FE_OFN1_scan_rst_sync1_mux_out),
	.SI(reg3[4]),
	.SE(n377),
	.Q(reg3[5]),
	.D(n278),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[3][0]  (
	.SI(reg2[7]),
	.SE(n377),
	.RN(rst),
	.Q(reg3[0]),
	.D(n273),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[3][1]  (
	.SI(reg3[0]),
	.SE(n380),
	.RN(rst),
	.Q(reg3[1]),
	.D(n274),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[3][4]  (
	.SI(reg3[3]),
	.SE(n379),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(reg3[4]),
	.D(n277),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[3][6]  (
	.SI(reg3[5]),
	.SE(n378),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(reg3[6]),
	.D(n279),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[3][3]  (
	.SI(reg3[2]),
	.SE(n377),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(reg3[3]),
	.D(n276),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[3][2]  (
	.SI(reg3[1]),
	.SE(n380),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(reg3[2]),
	.D(n275),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[3][7]  (
	.SI(reg3[6]),
	.SE(n379),
	.RN(FE_OFN1_scan_rst_sync1_mux_out),
	.Q(reg3[7]),
	.D(n280),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[2][4]  (
	.SI(test_si2),
	.SE(n378),
	.RN(rst),
	.Q(reg2[4]),
	.D(n285),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[2][2]  (
	.SI(reg2[1]),
	.SE(n377),
	.RN(rst),
	.Q(reg2[2]),
	.D(n283),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[2][5]  (
	.SI(reg2[4]),
	.SE(n379),
	.RN(rst),
	.Q(reg2[5]),
	.D(n286),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \reg_file_reg[2][6]  (
	.SI(reg2[5]),
	.SE(n378),
	.RN(rst),
	.Q(reg2[6]),
	.D(n287),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX1M \reg_file_reg[2][7]  (
	.SN(rst),
	.SI(reg2[6]),
	.SE(n380),
	.Q(reg2[7]),
	.D(n288),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3XLM U3 (
	.Y(n14),
	.C(N13),
	.B(n346),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3XLM U4 (
	.Y(n11),
	.C(N13),
	.B(n345),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4XLM U5 (
	.Y(N35),
	.S1(N12),
	.S0(N13),
	.D(n330),
	.C(n332),
	.B(n331),
	.A(n333), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4XLM U6 (
	.Y(N36),
	.S1(N12),
	.S0(N13),
	.D(n326),
	.C(n328),
	.B(n327),
	.A(n329), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4XLM U7 (
	.Y(N37),
	.S1(N12),
	.S0(N13),
	.D(n322),
	.C(n324),
	.B(n323),
	.A(n325), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4XLM U8 (
	.Y(N38),
	.S1(N12),
	.S0(N13),
	.D(n318),
	.C(n320),
	.B(n319),
	.A(n321), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3BX2M U9 (
	.Y(n29),
	.C(N13),
	.B(n345),
	.AN(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3BX2M U10 (
	.Y(n27),
	.C(n346),
	.B(N13),
	.AN(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U12 (
	.Y(n16),
	.B(N11),
	.A(n372), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U13 (
	.Y(n12),
	.B(n347),
	.A(n372), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U14 (
	.Y(n22),
	.B(N11),
	.A(N12), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U15 (
	.Y(n19),
	.B(N12),
	.A(n347), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U16 (
	.Y(n336),
	.A(n346), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U17 (
	.Y(n335),
	.A(n347), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U19 (
	.Y(n363),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U30 (
	.Y(n23),
	.B(rden),
	.AN(wren), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U32 (
	.Y(n26),
	.B(n12),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U34 (
	.Y(n28),
	.B(n12),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U36 (
	.Y(n32),
	.B(n16),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U38 (
	.Y(n33),
	.B(n16),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U40 (
	.Y(n34),
	.B(n19),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U42 (
	.Y(n35),
	.B(n19),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U44 (
	.Y(n36),
	.B(n22),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U46 (
	.Y(n37),
	.B(n22),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U47 (
	.Y(n15),
	.B(n11),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U48 (
	.Y(n17),
	.B(n14),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U49 (
	.Y(n18),
	.B(n11),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U50 (
	.Y(n20),
	.B(n14),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U51 (
	.Y(n21),
	.B(n11),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U52 (
	.Y(n24),
	.B(n14),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U53 (
	.Y(n13),
	.B(n12),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U54 (
	.Y(n2),
	.B(n12),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U55 (
	.Y(n364),
	.A(wrdata[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U56 (
	.Y(n1),
	.B(rden),
	.AN(wren), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U57 (
	.Y(n365),
	.A(wrdata[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U58 (
	.Y(n366),
	.A(wrdata[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U59 (
	.Y(n367),
	.A(wrdata[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U60 (
	.Y(n368),
	.A(wrdata[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U61 (
	.Y(n345),
	.A(n346), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U67 (
	.Y(n241),
	.B1(n26),
	.B0(n364),
	.A1N(n26),
	.A0N(\reg_file[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U68 (
	.Y(n242),
	.B1(n26),
	.B0(n365),
	.A1N(n26),
	.A0N(\reg_file[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U69 (
	.Y(n243),
	.B1(n26),
	.B0(n366),
	.A1N(n26),
	.A0N(\reg_file[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U70 (
	.Y(n244),
	.B1(n26),
	.B0(n367),
	.A1N(n26),
	.A0N(\reg_file[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U71 (
	.Y(n245),
	.B1(n26),
	.B0(n368),
	.A1N(n26),
	.A0N(\reg_file[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U72 (
	.Y(n246),
	.B1(n26),
	.B0(n369),
	.A1N(n26),
	.A0N(\reg_file[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U73 (
	.Y(n247),
	.B1(n26),
	.B0(n370),
	.A1N(n26),
	.A0N(\reg_file[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U74 (
	.Y(n248),
	.B1(n26),
	.B0(n371),
	.A1N(n26),
	.A0N(\reg_file[7][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U75 (
	.Y(n249),
	.B1(n28),
	.B0(n364),
	.A1N(n28),
	.A0N(\reg_file[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U76 (
	.Y(n250),
	.B1(n28),
	.B0(n365),
	.A1N(n28),
	.A0N(\reg_file[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U77 (
	.Y(n251),
	.B1(n28),
	.B0(n366),
	.A1N(n28),
	.A0N(\reg_file[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U78 (
	.Y(n252),
	.B1(n28),
	.B0(n367),
	.A1N(n28),
	.A0N(\reg_file[6][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U79 (
	.Y(n253),
	.B1(n28),
	.B0(n368),
	.A1N(n28),
	.A0N(\reg_file[6][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U80 (
	.Y(n254),
	.B1(n28),
	.B0(n369),
	.A1N(n28),
	.A0N(\reg_file[6][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U81 (
	.Y(n255),
	.B1(n28),
	.B0(n370),
	.A1N(n28),
	.A0N(\reg_file[6][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U82 (
	.Y(n256),
	.B1(n28),
	.B0(n371),
	.A1N(n28),
	.A0N(\reg_file[6][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U83 (
	.Y(n257),
	.B1(n32),
	.B0(n364),
	.A1N(n32),
	.A0N(\reg_file[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U84 (
	.Y(n258),
	.B1(n32),
	.B0(n365),
	.A1N(n32),
	.A0N(\reg_file[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U85 (
	.Y(n259),
	.B1(n32),
	.B0(n366),
	.A1N(n32),
	.A0N(\reg_file[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U86 (
	.Y(n260),
	.B1(n32),
	.B0(n367),
	.A1N(n32),
	.A0N(\reg_file[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U87 (
	.Y(n261),
	.B1(n32),
	.B0(n368),
	.A1N(n32),
	.A0N(\reg_file[5][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U88 (
	.Y(n262),
	.B1(n32),
	.B0(n369),
	.A1N(n32),
	.A0N(\reg_file[5][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U89 (
	.Y(n263),
	.B1(n32),
	.B0(n370),
	.A1N(n32),
	.A0N(\reg_file[5][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U90 (
	.Y(n264),
	.B1(n32),
	.B0(n371),
	.A1N(n32),
	.A0N(\reg_file[5][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U91 (
	.Y(n265),
	.B1(n33),
	.B0(n364),
	.A1N(n33),
	.A0N(\reg_file[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U92 (
	.Y(n266),
	.B1(n33),
	.B0(n365),
	.A1N(n33),
	.A0N(\reg_file[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U93 (
	.Y(n267),
	.B1(n33),
	.B0(n366),
	.A1N(n33),
	.A0N(\reg_file[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U94 (
	.Y(n268),
	.B1(n33),
	.B0(n367),
	.A1N(n33),
	.A0N(\reg_file[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U95 (
	.Y(n269),
	.B1(n33),
	.B0(n368),
	.A1N(n33),
	.A0N(\reg_file[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U96 (
	.Y(n270),
	.B1(n33),
	.B0(n369),
	.A1N(n33),
	.A0N(\reg_file[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U97 (
	.Y(n271),
	.B1(n33),
	.B0(n370),
	.A1N(n33),
	.A0N(\reg_file[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U98 (
	.Y(n272),
	.B1(n33),
	.B0(n371),
	.A1N(n33),
	.A0N(\reg_file[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U99 (
	.Y(n273),
	.B1(n34),
	.B0(n364),
	.A1N(n34),
	.A0N(reg3[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U100 (
	.Y(n274),
	.B1(n34),
	.B0(n365),
	.A1N(n34),
	.A0N(reg3[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U101 (
	.Y(n275),
	.B1(n34),
	.B0(n366),
	.A1N(n34),
	.A0N(reg3[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U102 (
	.Y(n276),
	.B1(n34),
	.B0(n367),
	.A1N(n34),
	.A0N(reg3[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U103 (
	.Y(n277),
	.B1(n34),
	.B0(n368),
	.A1N(n34),
	.A0N(reg3[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U104 (
	.Y(n279),
	.B1(n34),
	.B0(n370),
	.A1N(n34),
	.A0N(reg3[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U105 (
	.Y(n280),
	.B1(n34),
	.B0(n371),
	.A1N(n34),
	.A0N(reg3[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U106 (
	.Y(n282),
	.B1(n35),
	.B0(n365),
	.A1N(n35),
	.A0N(reg2[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U107 (
	.Y(n283),
	.B1(n35),
	.B0(n366),
	.A1N(n35),
	.A0N(reg2[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U108 (
	.Y(n284),
	.B1(n35),
	.B0(n367),
	.A1N(n35),
	.A0N(n384), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U109 (
	.Y(n285),
	.B1(n35),
	.B0(n368),
	.A1N(n35),
	.A0N(reg2[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U110 (
	.Y(n286),
	.B1(n35),
	.B0(n369),
	.A1N(n35),
	.A0N(reg2[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U111 (
	.Y(n287),
	.B1(n35),
	.B0(n370),
	.A1N(n35),
	.A0N(reg2[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U112 (
	.Y(n289),
	.B1(n36),
	.B0(n364),
	.A1N(n36),
	.A0N(reg1[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U113 (
	.Y(n290),
	.B1(n36),
	.B0(n365),
	.A1N(n36),
	.A0N(reg1[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U114 (
	.Y(n291),
	.B1(n36),
	.B0(n366),
	.A1N(n36),
	.A0N(reg1[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U115 (
	.Y(n292),
	.B1(n36),
	.B0(n367),
	.A1N(n36),
	.A0N(reg1[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U116 (
	.Y(n293),
	.B1(n36),
	.B0(n368),
	.A1N(n36),
	.A0N(reg1[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U117 (
	.Y(n294),
	.B1(n36),
	.B0(n369),
	.A1N(n36),
	.A0N(reg1[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U118 (
	.Y(n295),
	.B1(n36),
	.B0(n370),
	.A1N(n36),
	.A0N(reg1[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U119 (
	.Y(n296),
	.B1(n36),
	.B0(n371),
	.A1N(n36),
	.A0N(reg1[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U120 (
	.Y(n297),
	.B1(n37),
	.B0(n364),
	.A1N(n37),
	.A0N(reg0[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U121 (
	.Y(n298),
	.B1(n37),
	.B0(n365),
	.A1N(n37),
	.A0N(reg0[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U122 (
	.Y(n299),
	.B1(n37),
	.B0(n366),
	.A1N(n37),
	.A0N(reg0[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U123 (
	.Y(n300),
	.B1(n37),
	.B0(n367),
	.A1N(n37),
	.A0N(reg0[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U124 (
	.Y(n301),
	.B1(n37),
	.B0(n368),
	.A1N(n37),
	.A0N(reg0[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U125 (
	.Y(n302),
	.B1(n37),
	.B0(n369),
	.A1N(n37),
	.A0N(reg0[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U126 (
	.Y(n303),
	.B1(n37),
	.B0(n370),
	.A1N(n37),
	.A0N(reg0[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U127 (
	.Y(n304),
	.B1(n37),
	.B0(n371),
	.A1N(n37),
	.A0N(reg0[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U128 (
	.Y(n278),
	.B1(n34),
	.B0(n369),
	.A1N(n34),
	.A0N(reg3[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U129 (
	.Y(n281),
	.B1(n35),
	.B0(n364),
	.A1N(n35),
	.A0N(reg2[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U130 (
	.Y(n288),
	.B1(n35),
	.B0(n371),
	.A1N(n35),
	.A0N(reg2[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U131 (
	.Y(n369),
	.A(wrdata[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U132 (
	.Y(n370),
	.A(wrdata[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U133 (
	.Y(n371),
	.A(wrdata[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U134 (
	.Y(n209),
	.B1(n18),
	.B0(n364),
	.A1N(n18),
	.A0N(\reg_file[11][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U135 (
	.Y(n210),
	.B1(n18),
	.B0(n365),
	.A1N(n18),
	.A0N(\reg_file[11][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U136 (
	.Y(n211),
	.B1(n18),
	.B0(n366),
	.A1N(n18),
	.A0N(\reg_file[11][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U137 (
	.Y(n212),
	.B1(n18),
	.B0(n367),
	.A1N(n18),
	.A0N(\reg_file[11][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U138 (
	.Y(n213),
	.B1(n18),
	.B0(n368),
	.A1N(n18),
	.A0N(\reg_file[11][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U139 (
	.Y(n214),
	.B1(n18),
	.B0(n369),
	.A1N(n18),
	.A0N(\reg_file[11][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U140 (
	.Y(n215),
	.B1(n18),
	.B0(n370),
	.A1N(n18),
	.A0N(\reg_file[11][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U141 (
	.Y(n216),
	.B1(n18),
	.B0(n371),
	.A1N(n18),
	.A0N(\reg_file[11][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U142 (
	.Y(n217),
	.B1(n20),
	.B0(n364),
	.A1N(n20),
	.A0N(\reg_file[10][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U143 (
	.Y(n218),
	.B1(n20),
	.B0(n365),
	.A1N(n20),
	.A0N(\reg_file[10][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U144 (
	.Y(n219),
	.B1(n20),
	.B0(n366),
	.A1N(n20),
	.A0N(\reg_file[10][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U145 (
	.Y(n220),
	.B1(n20),
	.B0(n367),
	.A1N(n20),
	.A0N(\reg_file[10][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U146 (
	.Y(n221),
	.B1(n20),
	.B0(n368),
	.A1N(n20),
	.A0N(\reg_file[10][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U147 (
	.Y(n222),
	.B1(n20),
	.B0(n369),
	.A1N(n20),
	.A0N(\reg_file[10][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U148 (
	.Y(n223),
	.B1(n20),
	.B0(n370),
	.A1N(n20),
	.A0N(\reg_file[10][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U149 (
	.Y(n224),
	.B1(n20),
	.B0(n371),
	.A1N(n20),
	.A0N(\reg_file[10][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U150 (
	.Y(n225),
	.B1(n21),
	.B0(n364),
	.A1N(n21),
	.A0N(\reg_file[9][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U151 (
	.Y(n226),
	.B1(n21),
	.B0(n365),
	.A1N(n21),
	.A0N(\reg_file[9][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U152 (
	.Y(n227),
	.B1(n21),
	.B0(n366),
	.A1N(n21),
	.A0N(\reg_file[9][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U153 (
	.Y(n228),
	.B1(n21),
	.B0(n367),
	.A1N(n21),
	.A0N(\reg_file[9][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U154 (
	.Y(n229),
	.B1(n21),
	.B0(n368),
	.A1N(n21),
	.A0N(\reg_file[9][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U155 (
	.Y(n230),
	.B1(n21),
	.B0(n369),
	.A1N(n21),
	.A0N(\reg_file[9][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U156 (
	.Y(n231),
	.B1(n21),
	.B0(n370),
	.A1N(n21),
	.A0N(\reg_file[9][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U157 (
	.Y(n232),
	.B1(n21),
	.B0(n371),
	.A1N(n21),
	.A0N(\reg_file[9][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U158 (
	.Y(n233),
	.B1(n24),
	.B0(n364),
	.A1N(n24),
	.A0N(\reg_file[8][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U159 (
	.Y(n234),
	.B1(n24),
	.B0(n365),
	.A1N(n24),
	.A0N(\reg_file[8][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U160 (
	.Y(n235),
	.B1(n24),
	.B0(n366),
	.A1N(n24),
	.A0N(\reg_file[8][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U161 (
	.Y(n236),
	.B1(n24),
	.B0(n367),
	.A1N(n24),
	.A0N(\reg_file[8][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U162 (
	.Y(n237),
	.B1(n24),
	.B0(n368),
	.A1N(n24),
	.A0N(\reg_file[8][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U163 (
	.Y(n238),
	.B1(n24),
	.B0(n369),
	.A1N(n24),
	.A0N(\reg_file[8][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U164 (
	.Y(n239),
	.B1(n24),
	.B0(n370),
	.A1N(n24),
	.A0N(\reg_file[8][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U165 (
	.Y(n240),
	.B1(n24),
	.B0(n371),
	.A1N(n24),
	.A0N(\reg_file[8][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U166 (
	.Y(n193),
	.B1(n15),
	.B0(n364),
	.A1N(n15),
	.A0N(\reg_file[13][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U167 (
	.Y(n194),
	.B1(n15),
	.B0(n365),
	.A1N(n15),
	.A0N(\reg_file[13][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U168 (
	.Y(n195),
	.B1(n15),
	.B0(n366),
	.A1N(n15),
	.A0N(\reg_file[13][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U169 (
	.Y(n196),
	.B1(n15),
	.B0(n367),
	.A1N(n15),
	.A0N(\reg_file[13][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U170 (
	.Y(n197),
	.B1(n15),
	.B0(n368),
	.A1N(n15),
	.A0N(\reg_file[13][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U171 (
	.Y(n198),
	.B1(n15),
	.B0(n369),
	.A1N(n15),
	.A0N(\reg_file[13][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U172 (
	.Y(n199),
	.B1(n15),
	.B0(n370),
	.A1N(n15),
	.A0N(\reg_file[13][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U173 (
	.Y(n200),
	.B1(n15),
	.B0(n371),
	.A1N(n15),
	.A0N(\reg_file[13][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U174 (
	.Y(n201),
	.B1(n17),
	.B0(n364),
	.A1N(n17),
	.A0N(\reg_file[12][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U175 (
	.Y(n202),
	.B1(n17),
	.B0(n365),
	.A1N(n17),
	.A0N(\reg_file[12][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U176 (
	.Y(n203),
	.B1(n17),
	.B0(n366),
	.A1N(n17),
	.A0N(\reg_file[12][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U177 (
	.Y(n204),
	.B1(n17),
	.B0(n367),
	.A1N(n17),
	.A0N(\reg_file[12][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U315 (
	.Y(n205),
	.B1(n17),
	.B0(n368),
	.A1N(n17),
	.A0N(\reg_file[12][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U316 (
	.Y(n206),
	.B1(n17),
	.B0(n369),
	.A1N(n17),
	.A0N(n382), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U317 (
	.Y(n207),
	.B1(n17),
	.B0(n370),
	.A1N(n17),
	.A0N(\reg_file[12][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U318 (
	.Y(n208),
	.B1(n17),
	.B0(n371),
	.A1N(n17),
	.A0N(\reg_file[12][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U319 (
	.Y(n177),
	.B1(n364),
	.B0(n2),
	.A1N(n2),
	.A0N(\reg_file[15][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U320 (
	.Y(n178),
	.B1(n365),
	.B0(n2),
	.A1N(n2),
	.A0N(\reg_file[15][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U321 (
	.Y(n179),
	.B1(n366),
	.B0(n2),
	.A1N(n2),
	.A0N(\reg_file[15][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U322 (
	.Y(n180),
	.B1(n367),
	.B0(n2),
	.A1N(n2),
	.A0N(\reg_file[15][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U323 (
	.Y(n181),
	.B1(n368),
	.B0(n2),
	.A1N(n2),
	.A0N(\reg_file[15][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U324 (
	.Y(n182),
	.B1(n369),
	.B0(n2),
	.A1N(n2),
	.A0N(\reg_file[15][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U325 (
	.Y(n183),
	.B1(n370),
	.B0(n2),
	.A1N(n2),
	.A0N(\reg_file[15][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U326 (
	.Y(n184),
	.B1(n371),
	.B0(n2),
	.A1N(n2),
	.A0N(\reg_file[15][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U327 (
	.Y(n185),
	.B1(n13),
	.B0(n364),
	.A1N(n13),
	.A0N(\reg_file[14][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U328 (
	.Y(n186),
	.B1(n13),
	.B0(n365),
	.A1N(n13),
	.A0N(\reg_file[14][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U329 (
	.Y(n187),
	.B1(n13),
	.B0(n366),
	.A1N(n13),
	.A0N(\reg_file[14][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U330 (
	.Y(n188),
	.B1(n13),
	.B0(n367),
	.A1N(n13),
	.A0N(\reg_file[14][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U331 (
	.Y(n189),
	.B1(n13),
	.B0(n368),
	.A1N(n13),
	.A0N(\reg_file[14][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U332 (
	.Y(n190),
	.B1(n13),
	.B0(n369),
	.A1N(n13),
	.A0N(\reg_file[14][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U333 (
	.Y(n191),
	.B1(n13),
	.B0(n370),
	.A1N(n13),
	.A0N(\reg_file[14][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U334 (
	.Y(n192),
	.B1(n13),
	.B0(n371),
	.A1N(n13),
	.A0N(\reg_file[14][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U335 (
	.Y(n25),
	.S1(N11),
	.S0(n336),
	.D(reg3[1]),
	.C(reg2[1]),
	.B(reg1[1]),
	.A(reg0[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U336 (
	.Y(n6),
	.S1(N11),
	.S0(n345),
	.D(\reg_file[7][0] ),
	.C(\reg_file[6][0] ),
	.B(\reg_file[5][0] ),
	.A(\reg_file[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U337 (
	.Y(n10),
	.S1(N11),
	.S0(n336),
	.D(\reg_file[7][1] ),
	.C(\reg_file[6][1] ),
	.B(\reg_file[5][1] ),
	.A(\reg_file[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U338 (
	.Y(n38),
	.S1(n335),
	.S0(n336),
	.D(\reg_file[7][2] ),
	.C(\reg_file[6][2] ),
	.B(\reg_file[5][2] ),
	.A(\reg_file[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U339 (
	.Y(n316),
	.S1(n335),
	.S0(n336),
	.D(\reg_file[7][3] ),
	.C(\reg_file[6][3] ),
	.B(\reg_file[5][3] ),
	.A(\reg_file[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U340 (
	.Y(n320),
	.S1(n335),
	.S0(n336),
	.D(\reg_file[7][4] ),
	.C(\reg_file[6][4] ),
	.B(\reg_file[5][4] ),
	.A(\reg_file[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U341 (
	.Y(n324),
	.S1(N11),
	.S0(N10),
	.D(\reg_file[7][5] ),
	.C(\reg_file[6][5] ),
	.B(\reg_file[5][5] ),
	.A(\reg_file[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U342 (
	.Y(n328),
	.S1(N11),
	.S0(N10),
	.D(\reg_file[7][6] ),
	.C(\reg_file[6][6] ),
	.B(\reg_file[5][6] ),
	.A(\reg_file[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U343 (
	.Y(n332),
	.S1(N11),
	.S0(N10),
	.D(\reg_file[7][7] ),
	.C(\reg_file[6][7] ),
	.B(\reg_file[5][7] ),
	.A(\reg_file[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U344 (
	.Y(n4),
	.S1(N11),
	.S0(N10),
	.D(\reg_file[15][0] ),
	.C(\reg_file[14][0] ),
	.B(\reg_file[13][0] ),
	.A(\reg_file[12][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U345 (
	.Y(n30),
	.S1(n335),
	.S0(n336),
	.D(\reg_file[15][2] ),
	.C(\reg_file[14][2] ),
	.B(\reg_file[13][2] ),
	.A(\reg_file[12][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U346 (
	.Y(n314),
	.S1(n335),
	.S0(n336),
	.D(\reg_file[15][3] ),
	.C(\reg_file[14][3] ),
	.B(\reg_file[13][3] ),
	.A(\reg_file[12][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U347 (
	.Y(n318),
	.S1(n335),
	.S0(n336),
	.D(\reg_file[15][4] ),
	.C(\reg_file[14][4] ),
	.B(\reg_file[13][4] ),
	.A(\reg_file[12][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U348 (
	.Y(n322),
	.S1(N11),
	.S0(n345),
	.D(\reg_file[15][5] ),
	.C(\reg_file[14][5] ),
	.B(\reg_file[13][5] ),
	.A(n382), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U349 (
	.Y(n326),
	.S1(n335),
	.S0(N10),
	.D(\reg_file[15][6] ),
	.C(\reg_file[14][6] ),
	.B(\reg_file[13][6] ),
	.A(\reg_file[12][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U350 (
	.Y(n330),
	.S1(N11),
	.S0(N10),
	.D(\reg_file[15][7] ),
	.C(\reg_file[14][7] ),
	.B(\reg_file[13][7] ),
	.A(\reg_file[12][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U351 (
	.Y(n176),
	.B(n1),
	.AN(rddata_valid), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U352 (
	.Y(n305),
	.B1(n1),
	.B0(rddata[0]),
	.A1(n363),
	.A0(N42), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U353 (
	.Y(N42),
	.S1(N12),
	.S0(N13),
	.D(n4),
	.C(n6),
	.B(n5),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U354 (
	.Y(n7),
	.S1(N11),
	.S0(N10),
	.D(reg3[0]),
	.C(reg2[0]),
	.B(reg1[0]),
	.A(reg0[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U355 (
	.Y(n5),
	.S1(N11),
	.S0(N10),
	.D(\reg_file[11][0] ),
	.C(\reg_file[10][0] ),
	.B(\reg_file[9][0] ),
	.A(\reg_file[8][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U356 (
	.Y(n306),
	.B1(n1),
	.B0(rddata[1]),
	.A1(n363),
	.A0(N41), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U357 (
	.Y(N41),
	.S1(N12),
	.S0(N13),
	.D(n8),
	.C(n10),
	.B(n9),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U358 (
	.Y(n9),
	.S1(N11),
	.S0(N10),
	.D(\reg_file[11][1] ),
	.C(\reg_file[10][1] ),
	.B(\reg_file[9][1] ),
	.A(\reg_file[8][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U359 (
	.Y(n8),
	.S1(n335),
	.S0(n336),
	.D(\reg_file[15][1] ),
	.C(\reg_file[14][1] ),
	.B(\reg_file[13][1] ),
	.A(\reg_file[12][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U360 (
	.Y(n307),
	.B1(n1),
	.B0(rddata[2]),
	.A1(n363),
	.A0(N40), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U361 (
	.Y(N40),
	.S1(N12),
	.S0(N13),
	.D(n30),
	.C(n38),
	.B(n31),
	.A(n313), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U362 (
	.Y(n313),
	.S1(n335),
	.S0(n336),
	.D(reg3[2]),
	.C(reg2[2]),
	.B(reg1[2]),
	.A(reg0[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U363 (
	.Y(n31),
	.S1(n335),
	.S0(n336),
	.D(\reg_file[11][2] ),
	.C(\reg_file[10][2] ),
	.B(\reg_file[9][2] ),
	.A(\reg_file[8][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U364 (
	.Y(n308),
	.B1(n1),
	.B0(rddata[3]),
	.A1(n363),
	.A0(N39), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U365 (
	.Y(N39),
	.S1(N12),
	.S0(N13),
	.D(n314),
	.C(n316),
	.B(n315),
	.A(n317), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U366 (
	.Y(n317),
	.S1(n335),
	.S0(n336),
	.D(reg3[3]),
	.C(n384),
	.B(reg1[3]),
	.A(reg0[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U367 (
	.Y(n315),
	.S1(n335),
	.S0(n336),
	.D(\reg_file[11][3] ),
	.C(\reg_file[10][3] ),
	.B(\reg_file[9][3] ),
	.A(\reg_file[8][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U368 (
	.Y(n309),
	.B1(n1),
	.B0(rddata[4]),
	.A1(n363),
	.A0(N38), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U369 (
	.Y(n321),
	.S1(n335),
	.S0(N10),
	.D(reg3[4]),
	.C(reg2[4]),
	.B(reg1[4]),
	.A(reg0[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U370 (
	.Y(n319),
	.S1(n335),
	.S0(n336),
	.D(\reg_file[11][4] ),
	.C(\reg_file[10][4] ),
	.B(\reg_file[9][4] ),
	.A(\reg_file[8][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U371 (
	.Y(n310),
	.B1(n1),
	.B0(rddata[5]),
	.A1(n363),
	.A0(N37), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U372 (
	.Y(n325),
	.S1(N11),
	.S0(N10),
	.D(reg3[5]),
	.C(reg2[5]),
	.B(reg1[5]),
	.A(reg0[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U373 (
	.Y(n323),
	.S1(N11),
	.S0(N10),
	.D(\reg_file[11][5] ),
	.C(\reg_file[10][5] ),
	.B(\reg_file[9][5] ),
	.A(\reg_file[8][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U374 (
	.Y(n311),
	.B1(n1),
	.B0(rddata[6]),
	.A1(n363),
	.A0(N36), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U375 (
	.Y(n329),
	.S1(N11),
	.S0(n345),
	.D(reg3[6]),
	.C(reg2[6]),
	.B(reg1[6]),
	.A(reg0[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U376 (
	.Y(n327),
	.S1(N11),
	.S0(N10),
	.D(\reg_file[11][6] ),
	.C(\reg_file[10][6] ),
	.B(\reg_file[9][6] ),
	.A(\reg_file[8][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U377 (
	.Y(n312),
	.B1(n1),
	.B0(rddata[7]),
	.A1(n363),
	.A0(N35), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U378 (
	.Y(n333),
	.S1(N11),
	.S0(n345),
	.D(reg3[7]),
	.C(reg2[7]),
	.B(reg1[7]),
	.A(reg0[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U379 (
	.Y(n331),
	.S1(N11),
	.S0(N10),
	.D(\reg_file[11][7] ),
	.C(\reg_file[10][7] ),
	.B(\reg_file[9][7] ),
	.A(\reg_file[8][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U380 (
	.Y(n347),
	.A(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U381 (
	.Y(n346),
	.A(N10), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U382 (
	.Y(n372),
	.A(N12), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U383 (
	.Y(n377),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U384 (
	.Y(n378),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U385 (
	.Y(n379),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U386 (
	.Y(n380),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U387 (
	.Y(n381),
	.A(\reg_file[12][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U388 (
	.Y(n382),
	.A(n381), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U389 (
	.Y(n383),
	.A(reg2[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U390 (
	.Y(n384),
	.A(n383), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX4M \reg_file_reg[2][3]  (
	.SI(reg2[2]),
	.SE(n380),
	.RN(rst),
	.Q(FE_OFN11_SO_2_),
	.D(n284),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX4M \reg_file_reg[12][5]  (
	.SI(\reg_file[12][4] ),
	.SE(n377),
	.RN(FE_OFN2_scan_rst_sync1_mux_out),
	.Q(FE_OFN10_SO_1_),
	.D(n206),
	.CK(scan_clk_ref_clk_mux_out__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module bit16_alu_test_1 (
	a, 
	b, 
	alu_fun, 
	clk, 
	rst_n, 
	enable, 
	alu_out, 
	out_valid, 
	test_si, 
	test_se, 
	FE_OFN3_scan_rst_sync1_mux_out, 
	FE_OFN4_scan_rst_sync1_mux_out, 
	VDD, 
	VSS);
   input [7:0] a;
   input [7:0] b;
   input [3:0] alu_fun;
   input clk;
   input rst_n;
   input enable;
   output [15:0] alu_out;
   output out_valid;
   input test_si;
   input test_se;
   input FE_OFN3_scan_rst_sync1_mux_out;
   input FE_OFN4_scan_rst_sync1_mux_out;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_OFN7_n27;
   wire N92;
   wire N93;
   wire N94;
   wire N95;
   wire N96;
   wire N97;
   wire N98;
   wire N99;
   wire N100;
   wire N101;
   wire N102;
   wire N103;
   wire N104;
   wire N105;
   wire N106;
   wire N107;
   wire N108;
   wire N109;
   wire N110;
   wire N111;
   wire N112;
   wire N113;
   wire N114;
   wire N115;
   wire N116;
   wire N117;
   wire N118;
   wire N119;
   wire N120;
   wire N121;
   wire N122;
   wire N123;
   wire N124;
   wire N125;
   wire N126;
   wire N127;
   wire N128;
   wire N129;
   wire N130;
   wire N131;
   wire N132;
   wire N133;
   wire N158;
   wire N159;
   wire N160;
   wire N178;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n16;
   wire n18;
   wire n19;
   wire n21;
   wire n22;
   wire n24;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n33;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n58;
   wire n59;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n101;
   wire n102;
   wire n104;
   wire n105;
   wire n106;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n124;
   wire n126;
   wire n128;
   wire n130;
   wire n132;
   wire n134;
   wire n136;
   wire n138;
   wire n140;
   wire n142;
   wire n144;
   wire n146;
   wire n148;
   wire n150;
   wire n152;
   wire n154;
   wire n26;
   wire n32;
   wire n34;
   wire n40;
   wire n46;
   wire n47;
   wire n57;
   wire n60;
   wire n61;
   wire n68;
   wire n69;
   wire n76;
   wire n77;
   wire n84;
   wire n85;
   wire n93;
   wire n94;
   wire n100;
   wire n103;
   wire n107;
   wire n108;
   wire n109;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;

   // Module instantiations
   BUFX2M FE_OFC7_n27 (
	.Y(FE_OFN7_n27),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M out_valid_reg (
	.SI(alu_out[15]),
	.SE(test_se),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(out_valid),
	.D(N178),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \alu_out_reg[7]  (
	.SI(alu_out[6]),
	.SE(test_se),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(alu_out[7]),
	.D(n138),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \alu_out_reg[6]  (
	.SI(alu_out[5]),
	.SE(test_se),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(alu_out[6]),
	.D(n136),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \alu_out_reg[5]  (
	.SI(alu_out[4]),
	.SE(test_se),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(alu_out[5]),
	.D(n134),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \alu_out_reg[4]  (
	.SI(alu_out[3]),
	.SE(test_se),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(alu_out[4]),
	.D(n132),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \alu_out_reg[3]  (
	.SI(alu_out[2]),
	.SE(test_se),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(alu_out[3]),
	.D(n130),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX1M \alu_out_reg[2]  (
	.SI(alu_out[1]),
	.SE(test_se),
	.RN(rst_n),
	.Q(alu_out[2]),
	.D(n128),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX1M \alu_out_reg[1]  (
	.SI(alu_out[0]),
	.SE(test_se),
	.RN(rst_n),
	.Q(alu_out[1]),
	.D(n126),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX1M \alu_out_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(rst_n),
	.Q(alu_out[0]),
	.D(n124),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \alu_out_reg[15]  (
	.SI(alu_out[14]),
	.SE(test_se),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(alu_out[15]),
	.D(n154),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \alu_out_reg[14]  (
	.SI(alu_out[13]),
	.SE(test_se),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(alu_out[14]),
	.D(n152),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \alu_out_reg[13]  (
	.SI(alu_out[12]),
	.SE(test_se),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(alu_out[13]),
	.D(n150),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \alu_out_reg[12]  (
	.SI(alu_out[11]),
	.SE(test_se),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(alu_out[12]),
	.D(n148),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \alu_out_reg[11]  (
	.SI(alu_out[10]),
	.SE(test_se),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(alu_out[11]),
	.D(n146),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \alu_out_reg[10]  (
	.SI(alu_out[9]),
	.SE(test_se),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(alu_out[10]),
	.D(n144),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \alu_out_reg[9]  (
	.SI(alu_out[8]),
	.SE(test_se),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(alu_out[9]),
	.D(n142),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M \alu_out_reg[8]  (
	.SI(alu_out[7]),
	.SE(test_se),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(alu_out[8]),
	.D(n140),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U8 (
	.Y(n188),
	.A(enable), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U9 (
	.Y(n169),
	.A(n95), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U10 (
	.Y(n95),
	.B(n49),
	.A(n188), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U11 (
	.Y(n168),
	.A(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U12 (
	.Y(n166),
	.A(n44), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U13 (
	.Y(n49),
	.B1(n102),
	.B0(n171),
	.A1(n51),
	.A0(n175), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U14 (
	.Y(n90),
	.C(n176),
	.B(n188),
	.A(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U15 (
	.Y(n102),
	.B(n174),
	.A(n175), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U16 (
	.Y(n31),
	.B(n171),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U17 (
	.Y(n30),
	.B(n52),
	.A(enable), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U18 (
	.Y(n106),
	.B(n176),
	.A(n102), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U19 (
	.Y(n44),
	.B(n18),
	.A(n102), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U20 (
	.Y(n21),
	.B(n176),
	.A(n114), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U21 (
	.Y(n173),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U22 (
	.Y(n172),
	.A(FE_OFN7_n27), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U23 (
	.Y(n114),
	.B(n175),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U24 (
	.Y(n18),
	.C(n188),
	.B(alu_fun[0]),
	.A(n171), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U25 (
	.Y(n24),
	.D(n176),
	.C(n110),
	.B(alu_fun[3]),
	.A(enable), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U26 (
	.Y(n110),
	.B(alu_fun[1]),
	.A(alu_fun[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U27 (
	.Y(n101),
	.C(n188),
	.B(alu_fun[3]),
	.A(alu_fun[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U28 (
	.Y(n51),
	.C(n176),
	.B(alu_fun[2]),
	.A(n171), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U29 (
	.Y(n52),
	.B1(n43),
	.B0(alu_fun[3]),
	.A1N(n51),
	.A0N(n175), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U30 (
	.Y(n41),
	.B1(n187),
	.B0(n45),
	.A1(n44),
	.A0(n184), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U31 (
	.Y(n45),
	.B0(n168),
	.A1(n183),
	.A0(n173), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U32 (
	.Y(n33),
	.C(n176),
	.B(alu_fun[1]),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U33 (
	.Y(n29),
	.C(alu_fun[1]),
	.B(alu_fun[0]),
	.A(n101), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U34 (
	.Y(n43),
	.B(n175),
	.A(alu_fun[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U35 (
	.Y(n39),
	.B0(n172),
	.A1(n24),
	.A0(n183), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U36 (
	.Y(n171),
	.A(alu_fun[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U37 (
	.Y(n176),
	.A(alu_fun[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U38 (
	.Y(n175),
	.A(alu_fun[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U39 (
	.Y(n22),
	.B(alu_fun[0]),
	.A(n114), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U40 (
	.Y(n174),
	.A(alu_fun[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U41 (
	.Y(n14),
	.B(alu_fun[3]),
	.A(n90), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U42 (
	.Y(N178),
	.B(n188),
	.A(n122), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X2M U43 (
	.Y(n122),
	.D(n49),
	.C(alu_fun[2]),
	.B(n106),
	.A(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U45 (
	.Y(n27),
	.C(n106),
	.B(alu_fun[3]),
	.A(n188), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X2M U46 (
	.Y(n16),
	.D(alu_fun[1]),
	.C(n18),
	.B(n174),
	.A(N158), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U47 (
	.Y(n167),
	.A(n42), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M U48 (
	.Y(n42),
	.C(N160),
	.B(n18),
	.AN(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U49 (
	.Y(n126),
	.D(n38),
	.C(n37),
	.B(n36),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U50 (
	.Y(n38),
	.C0(n167),
	.B0(n41),
	.A1(n187),
	.A0(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U51 (
	.Y(n37),
	.C1(n21),
	.C0(N93),
	.B1(n14),
	.B0(a[2]),
	.A1(n22),
	.A0(N102), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U52 (
	.Y(n36),
	.C1(n29),
	.C0(N127),
	.B1(n48),
	.B0(enable),
	.A1(n183),
	.A0(FE_OFN7_n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U53 (
	.Y(n136),
	.D(n89),
	.C(n88),
	.B(n87),
	.A(n86), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U54 (
	.Y(n88),
	.C1(n163),
	.C0(n92),
	.B1(n22),
	.B0(N107),
	.A1(n91),
	.A0(b[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U55 (
	.Y(n89),
	.C1(n14),
	.C0(a[7]),
	.B1(n166),
	.B0(a[5]),
	.A1(n21),
	.A0(N98), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U56 (
	.Y(n87),
	.C1(n178),
	.C0(FE_OFN7_n27),
	.B1(n29),
	.B0(N132),
	.A1(n33),
	.A0(N116), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U57 (
	.Y(n111),
	.B0(n95),
	.A1(n22),
	.A0(N109), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U58 (
	.Y(n163),
	.A(b[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U59 (
	.Y(n105),
	.C0(FE_OFN7_n27),
	.B1(n177),
	.B0(n95),
	.A1(n173),
	.A0(a[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U60 (
	.Y(n104),
	.C0(n168),
	.B1(n170),
	.B0(a[7]),
	.A1(n177),
	.A0(n173), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U61 (
	.Y(n170),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U62 (
	.Y(n19),
	.C0(n172),
	.B1(n184),
	.B0(n24),
	.A1(n169),
	.A0(a[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U63 (
	.Y(n59),
	.C0(n172),
	.B1(n182),
	.B0(n24),
	.A1(n169),
	.A0(a[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U64 (
	.Y(n67),
	.C0(n172),
	.B1(n181),
	.B0(n24),
	.A1(n169),
	.A0(a[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U65 (
	.Y(n75),
	.C0(n172),
	.B1(n180),
	.B0(n24),
	.A1(n169),
	.A0(a[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U66 (
	.Y(n83),
	.C0(n172),
	.B1(n179),
	.B0(n24),
	.A1(n169),
	.A0(a[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U67 (
	.Y(n92),
	.C0(n172),
	.B1(n178),
	.B0(n24),
	.A1(n169),
	.A0(a[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U68 (
	.Y(n48),
	.B0(n50),
	.A2(a[1]),
	.A1(b[1]),
	.A0(n49), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI33X1M U69 (
	.Y(n50),
	.B2(b[1]),
	.B1(n52),
	.B0(a[1]),
	.A2(N159),
	.A1(alu_fun[1]),
	.A0(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U70 (
	.Y(n58),
	.C0(n31),
	.B1(n24),
	.B0(a[2]),
	.A1(n182),
	.A0(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U71 (
	.Y(n66),
	.C0(n31),
	.B1(n24),
	.B0(a[3]),
	.A1(n181),
	.A0(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U72 (
	.Y(n74),
	.C0(n31),
	.B1(n24),
	.B0(a[4]),
	.A1(n180),
	.A0(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U73 (
	.Y(n82),
	.C0(n31),
	.B1(n24),
	.B0(a[5]),
	.A1(n179),
	.A0(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U74 (
	.Y(n91),
	.C0(n31),
	.B1(n24),
	.B0(a[6]),
	.A1(n178),
	.A0(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U75 (
	.Y(n28),
	.C0(n31),
	.B1(n24),
	.B0(a[0]),
	.A1(n30),
	.A0(n184), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U76 (
	.Y(n164),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U77 (
	.Y(n165),
	.A(n76), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U78 (
	.Y(n177),
	.A(a[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U79 (
	.Y(n183),
	.A(a[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U80 (
	.Y(n184),
	.A(a[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U81 (
	.Y(n178),
	.A(a[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U82 (
	.Y(n181),
	.A(a[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U83 (
	.Y(n182),
	.A(a[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U84 (
	.Y(n180),
	.A(a[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U85 (
	.Y(n179),
	.A(a[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U86 (
	.Y(n187),
	.A(b[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U87 (
	.Y(n10),
	.C1(a[0]),
	.C0(n168),
	.B1(n33),
	.B0(N110),
	.A1(n188),
	.A0(alu_out[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U88 (
	.Y(n35),
	.C1(a[1]),
	.C0(n168),
	.B1(n33),
	.B0(N111),
	.A1(n188),
	.A0(alu_out[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U89 (
	.Y(n146),
	.B(n111),
	.A(n117), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U90 (
	.Y(n117),
	.B1(n188),
	.B0(alu_out[11]),
	.A1(n33),
	.A0(N121), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U91 (
	.Y(n150),
	.B(n111),
	.A(n119), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U92 (
	.Y(n119),
	.B1(n188),
	.B0(alu_out[13]),
	.A1(n33),
	.A0(N123), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U93 (
	.Y(n53),
	.B1(n188),
	.B0(alu_out[2]),
	.A1(n168),
	.A0(a[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U94 (
	.Y(n62),
	.B1(n188),
	.B0(alu_out[3]),
	.A1(n168),
	.A0(a[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U95 (
	.Y(n70),
	.B1(n188),
	.B0(alu_out[4]),
	.A1(n168),
	.A0(a[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U96 (
	.Y(n78),
	.B1(n188),
	.B0(alu_out[5]),
	.A1(n168),
	.A0(a[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U97 (
	.Y(n86),
	.B1(n188),
	.B0(alu_out[6]),
	.A1(n168),
	.A0(a[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U98 (
	.Y(n98),
	.B1(n188),
	.B0(alu_out[7]),
	.A1(n168),
	.A0(a[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U99 (
	.Y(n124),
	.D(n13),
	.C(n12),
	.B(n11),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U100 (
	.Y(n13),
	.C0(n16),
	.B0(n167),
	.A1(n14),
	.A0(a[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U101 (
	.Y(n12),
	.C1(n22),
	.C0(N101),
	.B1(n21),
	.B0(N92),
	.A1(n160),
	.A0(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X4M U102 (
	.Y(n11),
	.C1(n29),
	.C0(N126),
	.B1(n28),
	.B0(b[0]),
	.A1(n184),
	.A0(FE_OFN7_n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U103 (
	.Y(n128),
	.D(n56),
	.C(n55),
	.B(n54),
	.A(n53), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U104 (
	.Y(n55),
	.C1(n161),
	.C0(n59),
	.B1(n22),
	.B0(N103),
	.A1(n58),
	.A0(b[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U105 (
	.Y(n56),
	.C1(n14),
	.C0(a[3]),
	.B1(a[1]),
	.B0(n166),
	.A1(n21),
	.A0(N94), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U106 (
	.Y(n54),
	.C1(n182),
	.C0(FE_OFN7_n27),
	.B1(n29),
	.B0(N128),
	.A1(n33),
	.A0(N112), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U107 (
	.Y(n130),
	.D(n65),
	.C(n64),
	.B(n63),
	.A(n62), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U108 (
	.Y(n64),
	.C1(n162),
	.C0(n67),
	.B1(n22),
	.B0(N104),
	.A1(n66),
	.A0(b[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U109 (
	.Y(n65),
	.C1(n14),
	.C0(a[4]),
	.B1(n166),
	.B0(a[2]),
	.A1(n21),
	.A0(N95), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U110 (
	.Y(n63),
	.C1(n181),
	.C0(FE_OFN7_n27),
	.B1(n29),
	.B0(N129),
	.A1(n33),
	.A0(N113), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U111 (
	.Y(n132),
	.D(n73),
	.C(n72),
	.B(n71),
	.A(n70), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U112 (
	.Y(n72),
	.C1(n186),
	.C0(n75),
	.B1(n22),
	.B0(N105),
	.A1(n74),
	.A0(b[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U113 (
	.Y(n73),
	.C1(n14),
	.C0(a[5]),
	.B1(n166),
	.B0(a[3]),
	.A1(n21),
	.A0(N96), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U114 (
	.Y(n71),
	.C1(n180),
	.C0(FE_OFN7_n27),
	.B1(n29),
	.B0(N130),
	.A1(n33),
	.A0(N114), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U115 (
	.Y(n134),
	.D(n81),
	.C(n80),
	.B(n79),
	.A(n78), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U116 (
	.Y(n80),
	.C1(n185),
	.C0(n83),
	.B1(n22),
	.B0(N106),
	.A1(n82),
	.A0(b[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U117 (
	.Y(n81),
	.C1(n14),
	.C0(a[6]),
	.B1(n166),
	.B0(a[4]),
	.A1(n21),
	.A0(N97), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U118 (
	.Y(n79),
	.C1(n179),
	.C0(FE_OFN7_n27),
	.B1(n29),
	.B0(N131),
	.A1(n33),
	.A0(N115), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U119 (
	.Y(n142),
	.B(n111),
	.A(n115), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U120 (
	.Y(n115),
	.B1(n188),
	.B0(alu_out[9]),
	.A1(n33),
	.A0(N119), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U121 (
	.Y(n144),
	.B(n111),
	.A(n116), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U122 (
	.Y(n116),
	.B1(n188),
	.B0(alu_out[10]),
	.A1(n33),
	.A0(N120), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U123 (
	.Y(n148),
	.B(n111),
	.A(n118), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U124 (
	.Y(n118),
	.B1(n188),
	.B0(alu_out[12]),
	.A1(n33),
	.A0(N122), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U125 (
	.Y(n152),
	.B(n111),
	.A(n120), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U126 (
	.Y(n120),
	.B1(n188),
	.B0(alu_out[14]),
	.A1(n33),
	.A0(N124), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U127 (
	.Y(n154),
	.B(n111),
	.A(n121), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U128 (
	.Y(n121),
	.B1(n188),
	.B0(alu_out[15]),
	.A1(n33),
	.A0(N125), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U129 (
	.Y(n138),
	.D(n99),
	.C(n98),
	.B(n97),
	.AN(n96), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U130 (
	.Y(n96),
	.B1(n105),
	.B0(b[7]),
	.A1N(b[7]),
	.A0(n104), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U131 (
	.Y(n99),
	.C1(n177),
	.C0(FE_OFN7_n27),
	.B1(n29),
	.B0(N133),
	.A1(n33),
	.A0(N117), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U132 (
	.Y(n97),
	.C1(n21),
	.C0(N99),
	.B1(n166),
	.B0(a[6]),
	.A1(n22),
	.A0(N108), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B11X2M U133 (
	.Y(n140),
	.C0(n112),
	.B0(n111),
	.A1N(alu_out[8]),
	.A0(enable), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U134 (
	.Y(n112),
	.C0(n113),
	.B1(n21),
	.B0(N100),
	.A1(n33),
	.A0(N118), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U135 (
	.Y(n113),
	.C(n106),
	.B(n188),
	.A(n177), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U161 (
	.Y(n160),
	.A(b[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U162 (
	.Y(n161),
	.A(b[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U163 (
	.Y(n162),
	.A(b[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U164 (
	.Y(n186),
	.A(b[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U165 (
	.Y(n185),
	.A(b[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U166 (
	.Y(n156),
	.B(b[7]),
	.A(n177), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U167 (
	.Y(n93),
	.B(a[4]),
	.AN(b[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U168 (
	.Y(n46),
	.B(b[4]),
	.AN(a[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U169 (
	.Y(n100),
	.B(n46),
	.A(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U170 (
	.Y(n77),
	.B(a[3]),
	.A(n162), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U171 (
	.Y(n40),
	.B(a[2]),
	.A(n161), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U172 (
	.Y(n26),
	.B(a[0]),
	.A(n160), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U173 (
	.Y(n85),
	.B(n161),
	.A(a[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U174 (
	.Y(n68),
	.B(n85),
	.AN(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X1M U175 (
	.Y(n32),
	.B0(b[1]),
	.A1(n183),
	.A0(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X1M U176 (
	.Y(n34),
	.C0(n32),
	.B0(n68),
	.A1(n164),
	.A0(a[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U177 (
	.Y(n84),
	.B(n162),
	.A(a[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U178 (
	.Y(n47),
	.B0(n84),
	.A2(n34),
	.A1(n40),
	.A0(n77), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U179 (
	.Y(n108),
	.B(b[5]),
	.AN(a[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X1M U180 (
	.Y(n57),
	.C0(n108),
	.B0(n46),
	.A1(n47),
	.A0(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U181 (
	.Y(n94),
	.B(a[5]),
	.AN(b[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U182 (
	.Y(n107),
	.B(b[6]),
	.A(a[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U183 (
	.Y(n60),
	.B1(n178),
	.B0(b[6]),
	.A2(n107),
	.A1(n94),
	.A0(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U184 (
	.Y(n157),
	.B(n177),
	.A(b[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U185 (
	.Y(N160),
	.B0(n157),
	.A1(n60),
	.A0(n156), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U186 (
	.Y(n69),
	.B(n160),
	.A(a[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X1M U187 (
	.Y(n61),
	.B0(b[1]),
	.A1(n183),
	.A0(n69), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X1M U188 (
	.Y(n76),
	.C0(n61),
	.B0(n68),
	.A1(n183),
	.A0(n69), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X1M U189 (
	.Y(n103),
	.B0(n77),
	.A2(n84),
	.A1(n85),
	.A0(n165), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B11X1M U190 (
	.Y(n109),
	.C0(n93),
	.B0(n94),
	.A1N(n103),
	.A0(n100), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U191 (
	.Y(n158),
	.B1(n163),
	.B0(a[6]),
	.A2(n107),
	.A1(n108),
	.A0(n109), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2B1X1M U192 (
	.Y(n159),
	.B0(n156),
	.A1N(n158),
	.A0(n157), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U193 (
	.Y(N159),
	.A(n159), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U194 (
	.Y(N158),
	.B(N159),
	.A(N160), 
	.VDD(VDD), 
	.VSS(VSS));
   bit16_alu_DW_div_uns_0 div_30 (
	.a({ a[7],
		a[6],
		a[5],
		a[4],
		a[3],
		a[2],
		a[1],
		a[0] }),
	.b({ b[7],
		b[6],
		b[5],
		b[4],
		b[3],
		b[2],
		b[1],
		b[0] }),
	.quotient({ N133,
		N132,
		N131,
		N130,
		N129,
		N128,
		N127,
		N126 }),
	.n184(n184),
	.n183(n183),
	.n163(n163),
	.n182(n182), 
	.VDD(VDD), 
	.VSS(VSS));
   bit16_alu_DW01_sub_0 sub_24 (
	.A({ 1'b0,
		a[7],
		a[6],
		a[5],
		a[4],
		a[3],
		a[2],
		a[1],
		a[0] }),
	.B({ 1'b0,
		b[7],
		b[6],
		b[5],
		b[4],
		b[3],
		b[2],
		b[1],
		b[0] }),
	.CI(1'b0),
	.DIFF({ N109,
		N108,
		N107,
		N106,
		N105,
		N104,
		N103,
		N102,
		N101 }),
	.n160(n160),
	.n161(n161),
	.n162(n162),
	.n186(n186),
	.n185(n185),
	.n184(n184),
	.n187(n187),
	.n163(n163), 
	.VDD(VDD), 
	.VSS(VSS));
   bit16_alu_DW01_add_0 add_21 (
	.A({ 1'b0,
		a[7],
		a[6],
		a[5],
		a[4],
		a[3],
		a[2],
		a[1],
		a[0] }),
	.B({ 1'b0,
		b[7],
		b[6],
		b[5],
		b[4],
		b[3],
		b[2],
		b[1],
		b[0] }),
	.CI(1'b0),
	.SUM({ N100,
		N99,
		N98,
		N97,
		N96,
		N95,
		N94,
		N93,
		N92 }), 
	.VDD(VDD), 
	.VSS(VSS));
   bit16_alu_DW02_mult_0 mult_27 (
	.A({ a[7],
		a[6],
		a[5],
		a[4],
		a[3],
		a[2],
		a[1],
		a[0] }),
	.B({ b[7],
		b[6],
		b[5],
		b[4],
		b[3],
		b[2],
		b[1],
		b[0] }),
	.TC(1'b0),
	.PRODUCT({ N125,
		N124,
		N123,
		N122,
		N121,
		N120,
		N119,
		N118,
		N117,
		N116,
		N115,
		N114,
		N113,
		N112,
		N111,
		N110 }),
	.n160(n160),
	.n161(n161),
	.n162(n162),
	.n184(n184),
	.n183(n183),
	.n182(n182),
	.n181(n181),
	.n180(n180),
	.n179(n179),
	.n178(n178),
	.n177(n177),
	.n187(n187),
	.n163(n163),
	.n185(n185),
	.n186(n186), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module bit16_alu_DW_div_uns_0 (
	a, 
	b, 
	quotient, 
	remainder, 
	divide_by_0, 
	n184, 
	n183, 
	n163, 
	n182, 
	VDD, 
	VSS);
   input [7:0] a;
   input [7:0] b;
   output [7:0] quotient;
   output [7:0] remainder;
   output divide_by_0;
   input n184;
   input n183;
   input n163;
   input n182;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_RN_633_0;
   wire FE_RN_632_0;
   wire FE_RN_631_0;
   wire FE_RN_630_0;
   wire FE_RN_629_0;
   wire FE_RN_628_0;
   wire FE_RN_627_0;
   wire FE_RN_626_0;
   wire FE_RN_625_0;
   wire FE_RN_624_0;
   wire FE_RN_623_0;
   wire FE_RN_622_0;
   wire FE_RN_621_0;
   wire FE_RN_615_0;
   wire FE_RN_614_0;
   wire FE_RN_613_0;
   wire FE_RN_612_0;
   wire FE_RN_611_0;
   wire FE_RN_610_0;
   wire FE_RN_609_0;
   wire FE_RN_608_0;
   wire FE_RN_607_0;
   wire FE_RN_606_0;
   wire FE_RN_605_0;
   wire FE_RN_604_0;
   wire FE_RN_603_0;
   wire FE_RN_602_0;
   wire FE_RN_601_0;
   wire FE_RN_600_0;
   wire FE_RN_599_0;
   wire FE_RN_598_0;
   wire FE_RN_597_0;
   wire FE_RN_596_0;
   wire FE_RN_595_0;
   wire FE_RN_594_0;
   wire FE_RN_592_0;
   wire FE_RN_591_0;
   wire FE_RN_590_0;
   wire FE_RN_589_0;
   wire FE_RN_588_0;
   wire FE_RN_587_0;
   wire FE_RN_586_0;
   wire FE_RN_585_0;
   wire FE_RN_584_0;
   wire FE_RN_583_0;
   wire FE_RN_582_0;
   wire FE_RN_581_0;
   wire FE_RN_580_0;
   wire FE_RN_578_0;
   wire FE_RN_577_0;
   wire FE_RN_576_0;
   wire FE_RN_575_0;
   wire FE_RN_574_0;
   wire FE_RN_573_0;
   wire FE_RN_572_0;
   wire FE_RN_571_0;
   wire FE_RN_570_0;
   wire FE_RN_569_0;
   wire FE_RN_568_0;
   wire FE_RN_567_0;
   wire FE_RN_566_0;
   wire FE_RN_565_0;
   wire FE_RN_564_0;
   wire FE_RN_563_0;
   wire FE_RN_562_0;
   wire FE_RN_561_0;
   wire FE_RN_560_0;
   wire FE_RN_559_0;
   wire FE_RN_558_0;
   wire FE_RN_557_0;
   wire FE_RN_556_0;
   wire FE_RN_555_0;
   wire FE_RN_554_0;
   wire FE_RN_553_0;
   wire FE_RN_552_0;
   wire FE_RN_551_0;
   wire FE_RN_550_0;
   wire FE_RN_549_0;
   wire FE_RN_548_0;
   wire FE_RN_547_0;
   wire FE_RN_545_0;
   wire FE_RN_544_0;
   wire FE_RN_543_0;
   wire FE_RN_542_0;
   wire FE_RN_541_0;
   wire FE_RN_540_0;
   wire FE_RN_539_0;
   wire FE_RN_538_0;
   wire FE_RN_537_0;
   wire FE_RN_536_0;
   wire FE_RN_535_0;
   wire FE_RN_534_0;
   wire FE_RN_533_0;
   wire FE_RN_532_0;
   wire FE_RN_531_0;
   wire FE_RN_530_0;
   wire FE_RN_528_0;
   wire FE_RN_527_0;
   wire FE_RN_526_0;
   wire FE_RN_525_0;
   wire FE_RN_524_0;
   wire FE_RN_523_0;
   wire FE_RN_522_0;
   wire FE_RN_521_0;
   wire FE_RN_520_0;
   wire FE_RN_519_0;
   wire FE_RN_500_0;
   wire FE_RN_499_0;
   wire FE_RN_498_0;
   wire FE_RN_497_0;
   wire FE_RN_496_0;
   wire FE_RN_495_0;
   wire FE_RN_494_0;
   wire FE_RN_493_0;
   wire FE_RN_492_0;
   wire FE_RN_491_0;
   wire FE_RN_490_0;
   wire FE_RN_489_0;
   wire FE_RN_488_0;
   wire FE_RN_487_0;
   wire FE_RN_486_0;
   wire FE_RN_485_0;
   wire FE_RN_484_0;
   wire FE_RN_483_0;
   wire FE_RN_482_0;
   wire FE_RN_480_0;
   wire FE_RN_479_0;
   wire FE_RN_478_0;
   wire FE_RN_477_0;
   wire FE_RN_476_0;
   wire FE_RN_475_0;
   wire FE_RN_474_0;
   wire FE_RN_473_0;
   wire FE_RN_453_0;
   wire FE_RN_452_0;
   wire FE_RN_451_0;
   wire FE_RN_450_0;
   wire FE_RN_449_0;
   wire FE_RN_448_0;
   wire FE_RN_447_0;
   wire FE_RN_446_0;
   wire FE_RN_445_0;
   wire FE_RN_444_0;
   wire FE_RN_443_0;
   wire FE_RN_442_0;
   wire FE_RN_441_0;
   wire FE_RN_440_0;
   wire FE_RN_439_0;
   wire FE_RN_438_0;
   wire FE_RN_437_0;
   wire FE_RN_436_0;
   wire FE_RN_435_0;
   wire FE_RN_434_0;
   wire FE_RN_433_0;
   wire FE_RN_432_0;
   wire FE_RN_431_0;
   wire FE_RN_430_0;
   wire FE_RN_408_0;
   wire FE_RN_407_0;
   wire FE_RN_406_0;
   wire FE_RN_405_0;
   wire FE_RN_404_0;
   wire FE_RN_403_0;
   wire FE_RN_402_0;
   wire FE_RN_401_0;
   wire FE_RN_400_0;
   wire FE_RN_399_0;
   wire FE_RN_398_0;
   wire FE_RN_397_0;
   wire FE_RN_396_0;
   wire FE_RN_395_0;
   wire FE_RN_394_0;
   wire FE_RN_393_0;
   wire FE_RN_392_0;
   wire FE_RN_391_0;
   wire FE_RN_390_0;
   wire FE_RN_389_0;
   wire FE_RN_388_0;
   wire FE_RN_387_0;
   wire FE_RN_386_0;
   wire FE_RN_385_0;
   wire FE_RN_384_0;
   wire FE_RN_383_0;
   wire FE_RN_382_0;
   wire FE_RN_381_0;
   wire FE_RN_380_0;
   wire FE_RN_379_0;
   wire FE_RN_378_0;
   wire FE_RN_377_0;
   wire FE_RN_376_0;
   wire FE_RN_375_0;
   wire FE_RN_374_0;
   wire FE_RN_373_0;
   wire FE_RN_372_0;
   wire FE_RN_371_0;
   wire FE_RN_370_0;
   wire FE_RN_369_0;
   wire FE_RN_368_0;
   wire FE_RN_367_0;
   wire FE_RN_366_0;
   wire FE_RN_365_0;
   wire FE_RN_364_0;
   wire FE_RN_363_0;
   wire FE_RN_362_0;
   wire FE_RN_361_0;
   wire FE_RN_360_0;
   wire FE_RN_359_0;
   wire FE_RN_358_0;
   wire FE_RN_357_0;
   wire FE_RN_328_0;
   wire FE_RN_327_0;
   wire FE_RN_326_0;
   wire FE_RN_325_0;
   wire FE_RN_324_0;
   wire FE_RN_323_0;
   wire FE_RN_322_0;
   wire FE_RN_321_0;
   wire FE_RN_320_0;
   wire FE_RN_319_0;
   wire FE_RN_318_0;
   wire FE_RN_317_0;
   wire FE_RN_316_0;
   wire FE_RN_315_0;
   wire FE_RN_314_0;
   wire FE_RN_313_0;
   wire FE_RN_312_0;
   wire FE_RN_311_0;
   wire FE_RN_310_0;
   wire FE_RN_309_0;
   wire FE_RN_308_0;
   wire FE_RN_307_0;
   wire FE_RN_292_0;
   wire FE_RN_291_0;
   wire FE_RN_290_0;
   wire FE_RN_289_0;
   wire FE_RN_288_0;
   wire FE_RN_287_0;
   wire FE_RN_286_0;
   wire FE_RN_285_0;
   wire FE_RN_284_0;
   wire FE_RN_283_0;
   wire FE_RN_282_0;
   wire FE_RN_281_0;
   wire FE_RN_280_0;
   wire FE_RN_279_0;
   wire FE_RN_278_0;
   wire FE_RN_277_0;
   wire FE_RN_276_0;
   wire FE_RN_275_0;
   wire FE_RN_274_0;
   wire FE_RN_273_0;
   wire FE_RN_272_0;
   wire FE_RN_271_0;
   wire FE_RN_270_0;
   wire FE_RN_269_0;
   wire FE_RN_268_0;
   wire FE_RN_267_0;
   wire FE_RN_266_0;
   wire FE_RN_265_0;
   wire FE_RN_264_0;
   wire FE_RN_263_0;
   wire FE_RN_262_0;
   wire FE_RN_261_0;
   wire FE_RN_260_0;
   wire FE_RN_259_0;
   wire FE_RN_258_0;
   wire FE_RN_257_0;
   wire FE_RN_256_0;
   wire FE_RN_255_0;
   wire FE_RN_254_0;
   wire FE_RN_253_0;
   wire FE_RN_252_0;
   wire FE_RN_251_0;
   wire FE_RN_250_0;
   wire FE_RN_249_0;
   wire FE_RN_248_0;
   wire FE_RN_247_0;
   wire FE_RN_205_0;
   wire FE_RN_204_0;
   wire FE_RN_203_0;
   wire FE_RN_202_0;
   wire FE_RN_201_0;
   wire FE_RN_200_0;
   wire FE_RN_199_0;
   wire FE_RN_198_0;
   wire FE_RN_197_0;
   wire FE_RN_168_0;
   wire FE_RN_167_0;
   wire FE_RN_166_0;
   wire FE_RN_165_0;
   wire FE_RN_164_0;
   wire FE_RN_163_0;
   wire FE_RN_162_0;
   wire FE_RN_161_0;
   wire FE_RN_160_0;
   wire FE_RN_159_0;
   wire FE_RN_158_0;
   wire FE_RN_157_0;
   wire FE_RN_156_0;
   wire FE_RN_155_0;
   wire FE_RN_154_0;
   wire FE_RN_153_0;
   wire FE_RN_152_0;
   wire FE_RN_151_0;
   wire FE_RN_150_0;
   wire FE_RN_149_0;
   wire FE_RN_148_0;
   wire FE_RN_147_0;
   wire FE_RN_146_0;
   wire FE_RN_145_0;
   wire FE_RN_144_0;
   wire FE_RN_143_0;
   wire FE_RN_142_0;
   wire FE_RN_141_0;
   wire FE_RN_140_0;
   wire FE_RN_139_0;
   wire FE_RN_138_0;
   wire FE_RN_137_0;
   wire FE_RN_136_0;
   wire FE_RN_135_0;
   wire FE_RN_134_0;
   wire FE_RN_133_0;
   wire FE_RN_132_0;
   wire FE_RN_131_0;
   wire FE_RN_130_0;
   wire FE_RN_129_0;
   wire FE_RN_128_0;
   wire FE_RN_127_0;
   wire FE_RN_126_0;
   wire FE_RN_125_0;
   wire FE_RN_124_0;
   wire FE_RN_123_0;
   wire FE_RN_122_0;
   wire FE_RN_121_0;
   wire FE_RN_120_0;
   wire FE_RN_119_0;
   wire FE_RN_118_0;
   wire FE_RN_117_0;
   wire FE_RN_116_0;
   wire FE_RN_115_0;
   wire FE_RN_114_0;
   wire FE_RN_113_0;
   wire FE_RN_112_0;
   wire FE_RN_111_0;
   wire FE_RN_110_0;
   wire FE_RN_109_0;
   wire FE_RN_108_0;
   wire FE_RN_107_0;
   wire FE_RN_106_0;
   wire FE_RN_105_0;
   wire FE_RN_104_0;
   wire FE_RN_103_0;
   wire FE_RN_102_0;
   wire FE_RN_101_0;
   wire FE_RN_100_0;
   wire FE_RN_99_0;
   wire FE_RN_98_0;
   wire FE_RN_51_0;
   wire FE_RN_50_0;
   wire FE_RN_49_0;
   wire FE_RN_48_0;
   wire FE_RN_47_0;
   wire FE_RN_46_0;
   wire FE_RN_45_0;
   wire FE_RN_44_0;
   wire FE_RN_43_0;
   wire FE_RN_42_0;
   wire FE_RN_41_0;
   wire FE_RN_40_0;
   wire FE_RN_39_0;
   wire FE_RN_38_0;
   wire FE_RN_37_0;
   wire FE_RN_36_0;
   wire FE_RN_34_0;
   wire FE_RN_33_0;
   wire FE_RN_32_0;
   wire FE_RN_31_0;
   wire FE_RN_30_0;
   wire FE_RN_29_0;
   wire FE_RN_28_0;
   wire FE_RN_27_0;
   wire FE_RN_26_0;
   wire FE_RN_24_0;
   wire FE_RN_23_0;
   wire FE_RN_22_0;
   wire FE_RN_21_0;
   wire FE_RN_20_0;
   wire FE_RN_19_0;
   wire FE_RN_18_0;
   wire FE_RN_17_0;
   wire FE_RN_15_0;
   wire FE_RN_14_0;
   wire FE_RN_13_0;
   wire FE_RN_11_0;
   wire FE_RN_10_0;
   wire FE_RN_9_0;
   wire FE_RN_8_0;
   wire FE_RN_7_0;
   wire FE_RN_6_0;
   wire FE_RN_5_0;
   wire FE_RN_4_0;
   wire FE_RN_2_0;
   wire FE_RN_1_0;
   wire FE_RN_0_0;
   wire \u_div/SumTmp[1][0] ;
   wire \u_div/SumTmp[1][1] ;
   wire \u_div/SumTmp[1][2] ;
   wire \u_div/SumTmp[1][3] ;
   wire \u_div/SumTmp[1][4] ;
   wire \u_div/SumTmp[1][5] ;
   wire \u_div/SumTmp[1][6] ;
   wire \u_div/SumTmp[2][0] ;
   wire \u_div/SumTmp[2][1] ;
   wire \u_div/SumTmp[2][2] ;
   wire \u_div/SumTmp[2][3] ;
   wire \u_div/SumTmp[2][4] ;
   wire \u_div/SumTmp[2][5] ;
   wire \u_div/SumTmp[3][0] ;
   wire \u_div/SumTmp[3][1] ;
   wire \u_div/SumTmp[3][2] ;
   wire \u_div/SumTmp[3][3] ;
   wire \u_div/SumTmp[3][4] ;
   wire \u_div/SumTmp[4][0] ;
   wire \u_div/SumTmp[4][1] ;
   wire \u_div/SumTmp[4][2] ;
   wire \u_div/SumTmp[4][3] ;
   wire \u_div/SumTmp[5][0] ;
   wire \u_div/SumTmp[5][1] ;
   wire \u_div/SumTmp[5][2] ;
   wire \u_div/SumTmp[6][0] ;
   wire \u_div/SumTmp[7][0] ;
   wire \u_div/CryTmp[0][1] ;
   wire \u_div/CryTmp[0][2] ;
   wire \u_div/CryTmp[0][3] ;
   wire \u_div/CryTmp[0][4] ;
   wire \u_div/CryTmp[0][5] ;
   wire \u_div/CryTmp[0][6] ;
   wire \u_div/CryTmp[0][7] ;
   wire \u_div/CryTmp[1][1] ;
   wire \u_div/CryTmp[1][2] ;
   wire \u_div/CryTmp[2][1] ;
   wire \u_div/CryTmp[2][2] ;
   wire \u_div/CryTmp[2][3] ;
   wire \u_div/CryTmp[3][1] ;
   wire \u_div/CryTmp[3][2] ;
   wire \u_div/CryTmp[3][3] ;
   wire \u_div/CryTmp[4][1] ;
   wire \u_div/CryTmp[4][2] ;
   wire \u_div/CryTmp[4][3] ;
   wire \u_div/CryTmp[5][1] ;
   wire \u_div/CryTmp[5][2] ;
   wire \u_div/CryTmp[6][1] ;
   wire \u_div/CryTmp[7][1] ;
   wire \u_div/PartRem[1][1] ;
   wire \u_div/PartRem[1][2] ;
   wire \u_div/PartRem[1][3] ;
   wire \u_div/PartRem[1][4] ;
   wire \u_div/PartRem[1][5] ;
   wire \u_div/PartRem[1][6] ;
   wire \u_div/PartRem[1][7] ;
   wire \u_div/PartRem[2][1] ;
   wire \u_div/PartRem[2][2] ;
   wire \u_div/PartRem[2][3] ;
   wire \u_div/PartRem[2][4] ;
   wire \u_div/PartRem[2][5] ;
   wire \u_div/PartRem[2][6] ;
   wire \u_div/PartRem[3][1] ;
   wire \u_div/PartRem[3][2] ;
   wire \u_div/PartRem[3][3] ;
   wire \u_div/PartRem[3][4] ;
   wire \u_div/PartRem[3][5] ;
   wire \u_div/PartRem[4][1] ;
   wire \u_div/PartRem[4][2] ;
   wire \u_div/PartRem[4][3] ;
   wire \u_div/PartRem[4][4] ;
   wire \u_div/PartRem[5][1] ;
   wire \u_div/PartRem[5][2] ;
   wire \u_div/PartRem[5][3] ;
   wire \u_div/PartRem[6][1] ;
   wire \u_div/PartRem[6][2] ;
   wire \u_div/PartRem[7][1] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n12;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;

   // Module instantiations
   CLKAND2X12M FE_RC_738_0 (
	.Y(quotient[1]),
	.B(n12),
	.A(FE_RN_622_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_737_0 (
	.Y(FE_RN_633_0),
	.A(FE_RN_625_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_736_0 (
	.Y(FE_RN_632_0),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21BX4M FE_RC_735_0 (
	.Y(FE_RN_631_0),
	.B0N(FE_RN_632_0),
	.A1(FE_RN_633_0),
	.A0(FE_RN_627_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M FE_RC_734_0 (
	.Y(FE_RN_630_0),
	.B(FE_RN_580_0),
	.A(FE_RN_627_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_733_0 (
	.Y(FE_RN_629_0),
	.A(a[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21BX4M FE_RC_732_0 (
	.Y(FE_RN_628_0),
	.B0N(FE_RN_629_0),
	.A1(FE_RN_630_0),
	.A0(FE_RN_631_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_731_0 (
	.Y(FE_RN_627_0),
	.B(FE_RN_599_0),
	.A(FE_RN_597_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_730_0 (
	.Y(FE_RN_626_0),
	.A(FE_RN_627_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X3M FE_RC_729_0 (
	.Y(FE_RN_625_0),
	.B(FE_RN_586_0),
	.A(FE_RN_594_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_728_0 (
	.Y(FE_RN_624_0),
	.A(FE_RN_625_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_727_0 (
	.Y(FE_RN_623_0),
	.B(FE_RN_580_0),
	.A(FE_RN_624_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_726_0 (
	.Y(FE_RN_622_0),
	.B(FE_RN_626_0),
	.A(FE_RN_623_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M FE_RC_725_0 (
	.Y(FE_RN_621_0),
	.C(n12),
	.B(\u_div/SumTmp[1][0] ),
	.A(FE_RN_622_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_724_0 (
	.Y(\u_div/PartRem[1][1] ),
	.B(FE_RN_628_0),
	.A(FE_RN_621_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_717_0 (
	.Y(FE_RN_615_0),
	.A(FE_RN_589_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_716_0 (
	.Y(FE_RN_614_0),
	.B(FE_RN_615_0),
	.A(FE_RN_612_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_715_0 (
	.Y(FE_RN_613_0),
	.A(FE_RN_600_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_714_0 (
	.Y(FE_RN_612_0),
	.B(FE_RN_594_0),
	.A(FE_RN_613_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M FE_RC_713_0 (
	.Y(FE_RN_611_0),
	.C(FE_RN_586_0),
	.B(FE_RN_580_0),
	.A(FE_RN_612_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_712_0 (
	.Y(FE_RN_610_0),
	.A(FE_RN_580_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_711_0 (
	.Y(FE_RN_609_0),
	.A(FE_RN_603_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X3M FE_RC_710_0 (
	.Y(FE_RN_608_0),
	.C(FE_RN_589_0),
	.B(FE_RN_610_0),
	.A(FE_RN_609_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_709_0 (
	.Y(FE_RN_607_0),
	.A(FE_RN_586_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_708_0 (
	.Y(FE_RN_606_0),
	.A(n163), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_707_0 (
	.Y(FE_RN_605_0),
	.A(\u_div/PartRem[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_706_0 (
	.Y(FE_RN_604_0),
	.A(FE_RN_600_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M FE_RC_705_0 (
	.Y(FE_RN_603_0),
	.B0(FE_RN_604_0),
	.A1N(FE_RN_605_0),
	.A0N(FE_RN_606_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_704_0 (
	.Y(FE_RN_602_0),
	.A(FE_RN_603_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X3M FE_RC_703_0 (
	.Y(FE_RN_601_0),
	.C(FE_RN_589_0),
	.B(FE_RN_607_0),
	.A(FE_RN_602_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M FE_RC_702_0 (
	.Y(\u_div/SumTmp[1][6] ),
	.D(FE_RN_614_0),
	.C(FE_RN_611_0),
	.B(FE_RN_608_0),
	.A(FE_RN_601_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKAND2X6M FE_RC_701_0 (
	.Y(FE_RN_600_0),
	.B(n163),
	.A(\u_div/PartRem[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_700_0 (
	.Y(FE_RN_599_0),
	.A(FE_RN_600_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_699_0 (
	.Y(FE_RN_598_0),
	.A(FE_RN_589_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_698_0 (
	.Y(FE_RN_597_0),
	.B(FE_RN_598_0),
	.A(FE_RN_594_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_697_0 (
	.Y(FE_RN_596_0),
	.A(n163), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_696_0 (
	.Y(FE_RN_595_0),
	.A(\u_div/PartRem[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_695_0 (
	.Y(FE_RN_594_0),
	.B(FE_RN_596_0),
	.A(FE_RN_595_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M FE_RC_692_0 (
	.Y(FE_RN_592_0),
	.A(FE_RN_583_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X3M FE_RC_691_0 (
	.Y(FE_RN_525_0),
	.B(FE_RN_526_0),
	.A(FE_RN_592_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_690_0 (
	.Y(FE_RN_591_0),
	.B(n14),
	.A(\u_div/PartRem[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_689_0 (
	.Y(FE_RN_590_0),
	.B(FE_RN_591_0),
	.A(FE_RN_586_0), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M FE_RC_688_0 (
	.Y(\u_div/SumTmp[1][5] ),
	.B(FE_RN_590_0),
	.A(FE_RN_580_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_687_0 (
	.Y(FE_RN_589_0),
	.B(n14),
	.A(\u_div/PartRem[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_686_0 (
	.Y(FE_RN_588_0),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M FE_RC_685_0 (
	.Y(FE_RN_587_0),
	.A(\u_div/PartRem[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X3M FE_RC_684_0 (
	.Y(FE_RN_586_0),
	.B(FE_RN_588_0),
	.A(FE_RN_587_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_683_0 (
	.Y(FE_RN_585_0),
	.A(FE_RN_526_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_682_0 (
	.Y(FE_RN_584_0),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX4M FE_RC_681_0 (
	.Y(FE_RN_583_0),
	.B(FE_RN_584_0),
	.AN(\u_div/PartRem[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M FE_RC_680_0 (
	.Y(FE_RN_582_0),
	.D(FE_RN_547_0),
	.C(FE_RN_585_0),
	.B(FE_RN_550_0),
	.A(FE_RN_583_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X4M FE_RC_679_0 (
	.Y(FE_RN_581_0),
	.B(FE_RN_561_0),
	.A(FE_RN_557_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X3M FE_RC_678_0 (
	.Y(FE_RN_580_0),
	.C(FE_RN_555_0),
	.B(FE_RN_582_0),
	.A(FE_RN_581_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_675_0 (
	.Y(FE_RN_578_0),
	.A(FE_RN_554_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_674_0 (
	.Y(FE_RN_577_0),
	.B(\u_div/PartRem[2][1] ),
	.A(FE_RN_552_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX4M FE_RC_673_0 (
	.Y(\u_div/CryTmp[1][2] ),
	.B(FE_RN_577_0),
	.AN(FE_RN_578_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_672_0 (
	.Y(FE_RN_576_0),
	.A(FE_RN_568_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_671_0 (
	.Y(FE_RN_575_0),
	.A(FE_RN_554_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M FE_RC_670_0 (
	.Y(FE_RN_574_0),
	.B(\u_div/PartRem[2][1] ),
	.A(FE_RN_575_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_669_0 (
	.Y(FE_RN_573_0),
	.A(FE_RN_552_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M FE_RC_668_0 (
	.Y(FE_RN_572_0),
	.B(FE_RN_574_0),
	.A(FE_RN_573_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_667_0 (
	.Y(FE_RN_571_0),
	.B(FE_RN_525_0),
	.A(FE_RN_572_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_666_0 (
	.Y(FE_RN_570_0),
	.B(FE_RN_576_0),
	.A(FE_RN_571_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_665_0 (
	.Y(FE_RN_569_0),
	.A(FE_RN_550_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X3M FE_RC_664_0 (
	.Y(FE_RN_568_0),
	.B(FE_RN_530_0),
	.A(FE_RN_559_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2B1X2M FE_RC_663_0 (
	.Y(FE_RN_567_0),
	.B0(FE_RN_568_0),
	.A1N(FE_RN_569_0),
	.A0(FE_RN_525_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_662_0 (
	.Y(FE_RN_566_0),
	.B(n15),
	.A(\u_div/PartRem[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_661_0 (
	.Y(FE_RN_565_0),
	.B(FE_RN_547_0),
	.A(FE_RN_566_0), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M FE_RC_660_0 (
	.Y(\u_div/SumTmp[1][4] ),
	.S0(FE_RN_565_0),
	.B(FE_RN_567_0),
	.A(FE_RN_570_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M FE_RC_659_0 (
	.Y(FE_RN_564_0),
	.B1(\u_div/CryTmp[1][1] ),
	.B0(n18),
	.A1N(n18),
	.A0N(\u_div/CryTmp[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M FE_RC_658_0 (
	.Y(FE_RN_563_0),
	.B(FE_RN_554_0),
	.A(FE_RN_552_0), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X2M FE_RC_657_0 (
	.Y(\u_div/SumTmp[1][1] ),
	.S0(\u_div/PartRem[2][1] ),
	.B(FE_RN_563_0),
	.A(FE_RN_564_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_656_0 (
	.Y(FE_RN_562_0),
	.A(FE_RN_559_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_655_0 (
	.Y(FE_RN_561_0),
	.B(n15),
	.A(FE_RN_562_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_654_0 (
	.Y(FE_RN_560_0),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_653_0 (
	.Y(FE_RN_559_0),
	.B(FE_RN_519_0),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_652_0 (
	.Y(FE_RN_558_0),
	.B(FE_RN_560_0),
	.A(FE_RN_559_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_651_0 (
	.Y(FE_RN_557_0),
	.B(\u_div/PartRem[2][4] ),
	.A(FE_RN_558_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_650_0 (
	.Y(FE_RN_556_0),
	.A(FE_RN_530_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_649_0 (
	.Y(FE_RN_555_0),
	.B(FE_RN_556_0),
	.A(FE_RN_547_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_648_0 (
	.Y(FE_RN_554_0),
	.B(\u_div/CryTmp[1][1] ),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_647_0 (
	.Y(FE_RN_553_0),
	.A(FE_RN_554_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M FE_RC_646_0 (
	.Y(FE_RN_552_0),
	.B(\u_div/CryTmp[1][1] ),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_645_0 (
	.Y(FE_RN_551_0),
	.B(\u_div/PartRem[2][1] ),
	.A(FE_RN_552_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX4M FE_RC_644_0 (
	.Y(FE_RN_550_0),
	.B(FE_RN_551_0),
	.AN(FE_RN_553_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_643_0 (
	.Y(FE_RN_549_0),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_642_0 (
	.Y(FE_RN_548_0),
	.A(\u_div/PartRem[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_641_0 (
	.Y(FE_RN_547_0),
	.B(FE_RN_549_0),
	.A(FE_RN_548_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M FE_RC_638_0 (
	.Y(quotient[2]),
	.A(FE_RN_492_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_637_0 (
	.Y(FE_RN_545_0),
	.A(\u_div/SumTmp[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_636_0 (
	.Y(FE_RN_544_0),
	.A(\u_div/PartRem[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X2M FE_RC_635_0 (
	.Y(\u_div/PartRem[2][2] ),
	.S0(FE_RN_492_0),
	.B(FE_RN_544_0),
	.A(FE_RN_545_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_634_0 (
	.Y(FE_RN_543_0),
	.A(FE_RN_527_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_633_0 (
	.Y(FE_RN_542_0),
	.A(FE_RN_520_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2B1X4M FE_RC_632_0 (
	.Y(FE_RN_541_0),
	.B0(FE_RN_542_0),
	.A1N(FE_RN_543_0),
	.A0(\u_div/CryTmp[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X2M FE_RC_631_0 (
	.Y(FE_RN_540_0),
	.B(n16),
	.A(\u_div/PartRem[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B1X4M FE_RC_630_0 (
	.Y(FE_RN_539_0),
	.B0(FE_RN_527_0),
	.A1N(FE_RN_520_0),
	.A0(\u_div/CryTmp[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_629_0 (
	.Y(FE_RN_538_0),
	.B(FE_RN_540_0),
	.A(FE_RN_539_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X4M FE_RC_628_0 (
	.Y(\u_div/SumTmp[1][3] ),
	.B0(FE_RN_538_0),
	.A1(FE_RN_540_0),
	.A0(FE_RN_541_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_627_0 (
	.Y(FE_RN_537_0),
	.B(n17),
	.A(FE_RN_521_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M FE_RC_626_0 (
	.Y(FE_RN_536_0),
	.B0(FE_RN_537_0),
	.A1(n17),
	.A0(FE_RN_521_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_625_0 (
	.Y(FE_RN_535_0),
	.A(FE_RN_536_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_624_0 (
	.Y(FE_RN_534_0),
	.B(FE_RN_520_0),
	.A(FE_RN_527_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_623_0 (
	.Y(FE_RN_533_0),
	.B(\u_div/CryTmp[1][2] ),
	.A(FE_RN_534_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B1X2M FE_RC_622_0 (
	.Y(\u_div/SumTmp[1][2] ),
	.B0(FE_RN_533_0),
	.A1N(FE_RN_535_0),
	.A0(\u_div/CryTmp[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_621_0 (
	.Y(FE_RN_532_0),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X8M FE_RC_620_0 (
	.Y(FE_RN_531_0),
	.B(FE_RN_532_0),
	.A(FE_RN_520_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_619_0 (
	.Y(FE_RN_530_0),
	.B(\u_div/PartRem[2][3] ),
	.A(FE_RN_531_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_617_0 (
	.Y(FE_RN_528_0),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX8M FE_RC_616_0 (
	.Y(FE_RN_527_0),
	.B(FE_RN_528_0),
	.AN(FE_RN_521_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_615_0 (
	.Y(FE_RN_526_0),
	.A(FE_RN_527_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_613_0 (
	.Y(FE_RN_524_0),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_612_0 (
	.Y(FE_RN_523_0),
	.A(\u_div/SumTmp[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_611_0 (
	.Y(FE_RN_522_0),
	.A(\u_div/PartRem[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X6M FE_RC_610_0 (
	.Y(FE_RN_521_0),
	.S0(FE_RN_492_0),
	.B(FE_RN_522_0),
	.A(FE_RN_523_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX8M FE_RC_609_0 (
	.Y(FE_RN_520_0),
	.B(FE_RN_521_0),
	.AN(FE_RN_524_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_608_0 (
	.Y(FE_RN_519_0),
	.A(FE_RN_520_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M FE_RC_584_0 (
	.Y(FE_RN_482_0),
	.C(FE_RN_430_0),
	.B(\u_div/CryTmp[2][3] ),
	.A(FE_RN_433_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_582_0 (
	.Y(FE_RN_500_0),
	.A(\u_div/SumTmp[2][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_581_0 (
	.Y(FE_RN_499_0),
	.A(a[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_580_0 (
	.Y(FE_RN_498_0),
	.A(FE_RN_483_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_579_0 (
	.Y(FE_RN_497_0),
	.A(FE_RN_473_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X3M FE_RC_578_0 (
	.Y(FE_RN_496_0),
	.C(\u_div/CryTmp[2][3] ),
	.B(FE_RN_433_0),
	.A(FE_RN_430_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_577_0 (
	.Y(FE_RN_495_0),
	.B(FE_RN_435_0),
	.A(FE_RN_496_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_576_0 (
	.Y(FE_RN_494_0),
	.B(FE_RN_475_0),
	.A(FE_RN_495_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_575_0 (
	.Y(FE_RN_493_0),
	.B(FE_RN_497_0),
	.A(FE_RN_494_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_574_0 (
	.Y(FE_RN_492_0),
	.B(FE_RN_498_0),
	.A(FE_RN_493_0), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X4M FE_RC_573_0 (
	.Y(\u_div/PartRem[2][1] ),
	.S0(FE_RN_492_0),
	.B(FE_RN_499_0),
	.A(FE_RN_500_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_572_0 (
	.Y(FE_RN_491_0),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_571_0 (
	.Y(FE_RN_490_0),
	.A(\u_div/PartRem[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_570_0 (
	.Y(FE_RN_489_0),
	.A(FE_RN_479_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M FE_RC_569_0 (
	.Y(FE_RN_488_0),
	.B0(FE_RN_489_0),
	.A1N(FE_RN_490_0),
	.A0N(FE_RN_491_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_568_0 (
	.Y(FE_RN_487_0),
	.A(FE_RN_475_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X4M FE_RC_567_0 (
	.Y(FE_RN_486_0),
	.B(FE_RN_487_0),
	.A(FE_RN_479_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_566_0 (
	.Y(FE_RN_485_0),
	.A(FE_RN_438_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX4M FE_RC_565_0 (
	.Y(FE_RN_484_0),
	.C(FE_RN_435_0),
	.B(FE_RN_482_0),
	.AN(FE_RN_485_0), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X2M FE_RC_564_0 (
	.Y(\u_div/SumTmp[2][5] ),
	.S0(FE_RN_484_0),
	.B(FE_RN_486_0),
	.A(FE_RN_488_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_563_0 (
	.Y(FE_RN_483_0),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_560_0 (
	.Y(FE_RN_480_0),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX8M FE_RC_559_0 (
	.Y(FE_RN_479_0),
	.B(FE_RN_480_0),
	.AN(\u_div/PartRem[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_558_0 (
	.Y(FE_RN_478_0),
	.A(FE_RN_479_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_557_0 (
	.Y(FE_RN_477_0),
	.A(FE_RN_438_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_556_0 (
	.Y(FE_RN_476_0),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX8M FE_RC_555_0 (
	.Y(FE_RN_475_0),
	.B(FE_RN_476_0),
	.AN(\u_div/PartRem[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_554_0 (
	.Y(FE_RN_474_0),
	.B(FE_RN_477_0),
	.A(FE_RN_475_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_553_0 (
	.Y(FE_RN_473_0),
	.B(FE_RN_478_0),
	.A(FE_RN_474_0), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X2M FE_RC_530_0 (
	.Y(FE_RN_453_0),
	.B(n15),
	.A(\u_div/PartRem[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_529_0 (
	.Y(FE_RN_452_0),
	.A(\u_div/CryTmp[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_528_0 (
	.Y(FE_RN_451_0),
	.B(FE_RN_452_0),
	.A(FE_RN_437_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_527_0 (
	.Y(FE_RN_450_0),
	.B(FE_RN_433_0),
	.A(FE_RN_451_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_526_0 (
	.Y(FE_RN_449_0),
	.B(FE_RN_453_0),
	.A(FE_RN_450_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_525_0 (
	.Y(FE_RN_448_0),
	.A(FE_RN_437_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_524_0 (
	.Y(FE_RN_447_0),
	.B(FE_RN_448_0),
	.A(FE_RN_445_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_523_0 (
	.Y(FE_RN_446_0),
	.B(n15),
	.A(\u_div/PartRem[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_522_0 (
	.Y(FE_RN_445_0),
	.B(FE_RN_430_0),
	.A(FE_RN_446_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M FE_RC_521_0 (
	.Y(FE_RN_444_0),
	.C(\u_div/CryTmp[2][3] ),
	.B(FE_RN_433_0),
	.A(FE_RN_445_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M FE_RC_520_0 (
	.Y(\u_div/SumTmp[2][4] ),
	.C(FE_RN_449_0),
	.B(FE_RN_447_0),
	.A(FE_RN_444_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_519_0 (
	.Y(FE_RN_443_0),
	.A(\u_div/CryTmp[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X2M FE_RC_518_0 (
	.Y(FE_RN_442_0),
	.B(n16),
	.A(\u_div/PartRem[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_517_0 (
	.Y(FE_RN_441_0),
	.B(FE_RN_443_0),
	.A(FE_RN_442_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_516_0 (
	.Y(FE_RN_440_0),
	.B(FE_RN_437_0),
	.A(FE_RN_433_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_515_0 (
	.Y(FE_RN_439_0),
	.B(\u_div/CryTmp[2][3] ),
	.A(FE_RN_440_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_514_0 (
	.Y(\u_div/SumTmp[2][3] ),
	.B(FE_RN_441_0),
	.A(FE_RN_439_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_513_0 (
	.Y(FE_RN_438_0),
	.B(n15),
	.A(\u_div/PartRem[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_512_0 (
	.Y(FE_RN_437_0),
	.B(n16),
	.A(\u_div/PartRem[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_511_0 (
	.Y(FE_RN_436_0),
	.A(FE_RN_437_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_510_0 (
	.Y(FE_RN_435_0),
	.B(FE_RN_436_0),
	.A(FE_RN_430_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_509_0 (
	.Y(FE_RN_434_0),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX8M FE_RC_508_0 (
	.Y(FE_RN_433_0),
	.B(FE_RN_434_0),
	.AN(\u_div/PartRem[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_507_0 (
	.Y(FE_RN_432_0),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_506_0 (
	.Y(FE_RN_431_0),
	.A(\u_div/PartRem[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_505_0 (
	.Y(FE_RN_430_0),
	.B(FE_RN_432_0),
	.A(FE_RN_431_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_479_0 (
	.Y(FE_RN_408_0),
	.A(FE_RN_383_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X12M FE_RC_478_0 (
	.Y(quotient[3]),
	.B(FE_RN_408_0),
	.A(FE_RN_387_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X3M FE_RC_477_0 (
	.Y(FE_RN_407_0),
	.B(FE_RN_387_0),
	.A(FE_RN_382_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_476_0 (
	.Y(FE_RN_406_0),
	.B(\u_div/PartRem[4][1] ),
	.A(FE_RN_404_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X3M FE_RC_475_0 (
	.Y(\u_div/PartRem[3][2] ),
	.B(FE_RN_407_0),
	.A(FE_RN_406_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_474_0 (
	.Y(FE_RN_405_0),
	.A(FE_RN_383_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X6M FE_RC_473_0 (
	.Y(FE_RN_404_0),
	.B(FE_RN_405_0),
	.A(FE_RN_387_0), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X4M FE_RC_472_0 (
	.Y(FE_RN_403_0),
	.B(\u_div/PartRem[4][1] ),
	.A(FE_RN_399_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_471_0 (
	.Y(FE_RN_402_0),
	.B(FE_RN_404_0),
	.A(FE_RN_403_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_470_0 (
	.Y(FE_RN_401_0),
	.A(FE_RN_383_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_469_0 (
	.Y(FE_RN_400_0),
	.A(\u_div/CryTmp[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X4M FE_RC_468_0 (
	.Y(FE_RN_399_0),
	.S0(n17),
	.B(FE_RN_400_0),
	.A(\u_div/CryTmp[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X4M FE_RC_467_0 (
	.Y(FE_RN_398_0),
	.B(\u_div/SumTmp[3][1] ),
	.A(FE_RN_399_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M FE_RC_466_0 (
	.Y(FE_RN_397_0),
	.C(FE_RN_401_0),
	.B(FE_RN_387_0),
	.A(FE_RN_398_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_465_0 (
	.Y(\u_div/SumTmp[2][2] ),
	.B(FE_RN_402_0),
	.A(FE_RN_397_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_464_0 (
	.Y(FE_RN_396_0),
	.A(FE_RN_307_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_463_0 (
	.Y(FE_RN_395_0),
	.A(\u_div/PartRem[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X4M FE_RC_462_0 (
	.Y(FE_RN_394_0),
	.B(FE_RN_395_0),
	.A(FE_RN_387_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_461_0 (
	.Y(FE_RN_393_0),
	.B(\u_div/PartRem[4][1] ),
	.A(FE_RN_383_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_460_0 (
	.Y(FE_RN_392_0),
	.B(FE_RN_386_0),
	.A(FE_RN_382_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_459_0 (
	.Y(FE_RN_391_0),
	.B(FE_RN_393_0),
	.A(FE_RN_392_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X4M FE_RC_458_0 (
	.Y(FE_RN_390_0),
	.C0(FE_RN_391_0),
	.B0(FE_RN_394_0),
	.A1(FE_RN_396_0),
	.A0(FE_RN_382_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_457_0 (
	.Y(FE_RN_389_0),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_456_0 (
	.Y(FE_RN_388_0),
	.A(FE_RN_386_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X6M FE_RC_455_0 (
	.Y(FE_RN_387_0),
	.B(FE_RN_307_0),
	.A(FE_RN_388_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X5M FE_RC_454_0 (
	.Y(FE_RN_386_0),
	.B(FE_RN_316_0),
	.A(FE_RN_312_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21X2M FE_RC_453_0 (
	.Y(FE_RN_385_0),
	.B0(n17),
	.A1(\u_div/PartRem[4][1] ),
	.A0(FE_RN_383_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X1M FE_RC_452_0 (
	.Y(FE_RN_384_0),
	.B0(FE_RN_385_0),
	.A1(FE_RN_386_0),
	.A0(FE_RN_382_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_451_0 (
	.Y(FE_RN_383_0),
	.B(n14),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M FE_RC_450_0 (
	.Y(FE_RN_382_0),
	.B(FE_RN_383_0),
	.AN(\u_div/SumTmp[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M FE_RC_449_0 (
	.Y(FE_RN_381_0),
	.B(FE_RN_382_0),
	.AN(FE_RN_307_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B11X4M FE_RC_448_0 (
	.Y(FE_RN_380_0),
	.C0(FE_RN_381_0),
	.B0(FE_RN_384_0),
	.A1N(\u_div/PartRem[4][1] ),
	.A0(FE_RN_387_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X3M FE_RC_447_0 (
	.Y(FE_RN_379_0),
	.B(\u_div/CryTmp[2][2] ),
	.A(FE_RN_380_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X4M FE_RC_446_0 (
	.Y(\u_div/CryTmp[2][3] ),
	.B0(FE_RN_379_0),
	.A1(FE_RN_389_0),
	.A0(FE_RN_390_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_445_0 (
	.Y(FE_RN_378_0),
	.A(a[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_444_0 (
	.Y(FE_RN_377_0),
	.A(\u_div/SumTmp[3][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X6M FE_RC_443_0 (
	.Y(\u_div/PartRem[3][1] ),
	.S0(quotient[3]),
	.B(FE_RN_377_0),
	.A(FE_RN_378_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_442_0 (
	.Y(FE_RN_376_0),
	.A(FE_RN_372_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_441_0 (
	.Y(FE_RN_375_0),
	.A(a[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_440_0 (
	.Y(FE_RN_374_0),
	.A(a[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_439_0 (
	.Y(FE_RN_373_0),
	.B(n18),
	.A(FE_RN_374_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X4M FE_RC_438_0 (
	.Y(FE_RN_372_0),
	.B0(FE_RN_373_0),
	.A1(n18),
	.A0(FE_RN_375_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_437_0 (
	.Y(FE_RN_371_0),
	.A(FE_RN_372_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_436_0 (
	.Y(FE_RN_370_0),
	.B(\u_div/CryTmp[2][1] ),
	.A(FE_RN_371_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M FE_RC_435_0 (
	.Y(FE_RN_369_0),
	.B0(FE_RN_370_0),
	.A1(\u_div/CryTmp[2][1] ),
	.A0(FE_RN_376_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_434_0 (
	.Y(FE_RN_368_0),
	.A(\u_div/CryTmp[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_433_0 (
	.Y(FE_RN_367_0),
	.A(\u_div/CryTmp[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X4M FE_RC_432_0 (
	.Y(FE_RN_366_0),
	.B(n18),
	.A(\u_div/SumTmp[3][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_431_0 (
	.Y(FE_RN_365_0),
	.B(FE_RN_367_0),
	.A(FE_RN_366_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X4M FE_RC_430_0 (
	.Y(FE_RN_364_0),
	.B0(FE_RN_365_0),
	.A1(FE_RN_368_0),
	.A0(FE_RN_366_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_429_0 (
	.Y(FE_RN_363_0),
	.B(quotient[3]),
	.A(FE_RN_364_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B1X4M FE_RC_428_0 (
	.Y(\u_div/SumTmp[2][1] ),
	.B0(FE_RN_363_0),
	.A1N(FE_RN_369_0),
	.A0(quotient[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X4M FE_RC_427_0 (
	.Y(FE_RN_362_0),
	.B(a[3]),
	.A(FE_RN_360_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_426_0 (
	.Y(FE_RN_361_0),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX8M FE_RC_425_0 (
	.Y(FE_RN_360_0),
	.B(FE_RN_361_0),
	.AN(\u_div/CryTmp[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X4M FE_RC_424_0 (
	.Y(FE_RN_359_0),
	.B(\u_div/SumTmp[3][0] ),
	.A(FE_RN_360_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X8M FE_RC_423_0 (
	.Y(FE_RN_358_0),
	.B(quotient[3]),
	.A(FE_RN_359_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_422_0 (
	.Y(FE_RN_357_0),
	.B(\u_div/CryTmp[2][1] ),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B11X4M FE_RC_421_0 (
	.Y(\u_div/CryTmp[2][2] ),
	.C0(FE_RN_357_0),
	.B0(FE_RN_358_0),
	.A1N(FE_RN_362_0),
	.A0(quotient[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_386_0 (
	.Y(FE_RN_328_0),
	.A(\u_div/PartRem[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M FE_RC_385_0 (
	.Y(\u_div/PartRem[4][3] ),
	.B1(quotient[4]),
	.B0(FE_RN_328_0),
	.A1N(\u_div/SumTmp[4][2] ),
	.A0N(quotient[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_384_0 (
	.Y(FE_RN_327_0),
	.A(\u_div/CryTmp[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_383_0 (
	.Y(FE_RN_326_0),
	.A(FE_RN_314_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2B1X8M FE_RC_382_0 (
	.Y(FE_RN_325_0),
	.B0(FE_RN_326_0),
	.A1N(FE_RN_327_0),
	.A0(FE_RN_308_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_381_0 (
	.Y(FE_RN_324_0),
	.A(FE_RN_308_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2B1X2M FE_RC_380_0 (
	.Y(FE_RN_323_0),
	.B0(FE_RN_324_0),
	.A1N(\u_div/CryTmp[3][3] ),
	.A0(FE_RN_314_0), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X4M FE_RC_379_0 (
	.Y(FE_RN_322_0),
	.B(n15),
	.A(\u_div/PartRem[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X2M FE_RC_378_0 (
	.Y(\u_div/SumTmp[3][4] ),
	.S0(FE_RN_322_0),
	.B(FE_RN_323_0),
	.A(FE_RN_325_0), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M FE_RC_377_0 (
	.Y(FE_RN_321_0),
	.B(n16),
	.A(FE_RN_310_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_376_0 (
	.Y(FE_RN_320_0),
	.B(FE_RN_314_0),
	.A(FE_RN_308_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_375_0 (
	.Y(FE_RN_319_0),
	.B(\u_div/CryTmp[3][3] ),
	.A(FE_RN_320_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X4M FE_RC_374_0 (
	.Y(\u_div/SumTmp[3][3] ),
	.B0(FE_RN_319_0),
	.A1(\u_div/CryTmp[3][3] ),
	.A0(FE_RN_321_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_373_0 (
	.Y(FE_RN_318_0),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_372_0 (
	.Y(FE_RN_317_0),
	.B(FE_RN_318_0),
	.A(FE_RN_314_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_371_0 (
	.Y(FE_RN_316_0),
	.B(\u_div/PartRem[4][4] ),
	.A(FE_RN_317_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_370_0 (
	.Y(FE_RN_315_0),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X8M FE_RC_369_0 (
	.Y(FE_RN_314_0),
	.B(n16),
	.A(FE_RN_310_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_368_0 (
	.Y(FE_RN_313_0),
	.A(FE_RN_314_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M FE_RC_367_0 (
	.Y(FE_RN_312_0),
	.B(FE_RN_313_0),
	.AN(FE_RN_315_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_366_0 (
	.Y(FE_RN_311_0),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M FE_RC_365_0 (
	.Y(FE_RN_310_0),
	.S0(quotient[4]),
	.B(\u_div/SumTmp[4][2] ),
	.A(\u_div/PartRem[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_364_0 (
	.Y(FE_RN_309_0),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX8M FE_RC_363_0 (
	.Y(FE_RN_308_0),
	.B(FE_RN_309_0),
	.AN(FE_RN_310_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B11X4M FE_RC_362_0 (
	.Y(FE_RN_307_0),
	.C0(\u_div/CryTmp[3][3] ),
	.B0(FE_RN_308_0),
	.A1N(FE_RN_311_0),
	.A0(\u_div/PartRem[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X8M FE_RC_342_0 (
	.Y(quotient[4]),
	.B(FE_RN_197_0),
	.A(FE_RN_200_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_341_0 (
	.Y(FE_RN_292_0),
	.B(\u_div/SumTmp[4][1] ),
	.A(FE_RN_279_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX8M FE_RC_340_0 (
	.Y(\u_div/PartRem[4][2] ),
	.B(FE_RN_292_0),
	.AN(FE_RN_278_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_339_0 (
	.Y(FE_RN_291_0),
	.A(\u_div/CryTmp[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_338_0 (
	.Y(FE_RN_290_0),
	.A(\u_div/PartRem[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_337_0 (
	.Y(FE_RN_289_0),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M FE_RC_336_0 (
	.Y(FE_RN_288_0),
	.B1(\u_div/PartRem[5][1] ),
	.B0(FE_RN_289_0),
	.A1(n17),
	.A0(FE_RN_290_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_335_0 (
	.Y(FE_RN_287_0),
	.A(\u_div/SumTmp[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_334_0 (
	.Y(FE_RN_286_0),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M FE_RC_333_0 (
	.Y(FE_RN_285_0),
	.B1(\u_div/SumTmp[4][1] ),
	.B0(FE_RN_286_0),
	.A1(n17),
	.A0(FE_RN_287_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_332_0 (
	.Y(FE_RN_284_0),
	.B(FE_RN_285_0),
	.A(FE_RN_279_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X4M FE_RC_331_0 (
	.Y(FE_RN_283_0),
	.B0(FE_RN_284_0),
	.A1(FE_RN_288_0),
	.A0(FE_RN_279_0), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X4M FE_RC_330_0 (
	.Y(\u_div/SumTmp[3][2] ),
	.S0(FE_RN_283_0),
	.B(\u_div/CryTmp[3][2] ),
	.A(FE_RN_291_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_329_0 (
	.Y(FE_RN_282_0),
	.B(\u_div/SumTmp[4][1] ),
	.A(FE_RN_279_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B1X8M FE_RC_328_0 (
	.Y(FE_RN_281_0),
	.B0(n17),
	.A1N(FE_RN_282_0),
	.A0(FE_RN_278_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_327_0 (
	.Y(FE_RN_280_0),
	.A(\u_div/PartRem[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_326_0 (
	.Y(FE_RN_279_0),
	.B(FE_RN_200_0),
	.A(FE_RN_197_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X8M FE_RC_325_0 (
	.Y(FE_RN_278_0),
	.B(FE_RN_280_0),
	.A(FE_RN_279_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_324_0 (
	.Y(FE_RN_277_0),
	.A(\u_div/SumTmp[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_323_0 (
	.Y(FE_RN_276_0),
	.A(\u_div/SumTmp[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_322_0 (
	.Y(FE_RN_275_0),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M FE_RC_321_0 (
	.Y(FE_RN_274_0),
	.B0(FE_RN_275_0),
	.A1(FE_RN_200_0),
	.A0(FE_RN_276_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X4M FE_RC_320_0 (
	.Y(FE_RN_273_0),
	.B0(FE_RN_274_0),
	.A1N(FE_RN_197_0),
	.A0N(FE_RN_277_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX8M FE_RC_319_0 (
	.Y(FE_RN_272_0),
	.B(FE_RN_273_0),
	.AN(FE_RN_278_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_318_0 (
	.Y(FE_RN_271_0),
	.B(\u_div/CryTmp[3][2] ),
	.A(FE_RN_272_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_317_0 (
	.Y(\u_div/CryTmp[3][3] ),
	.B(FE_RN_281_0),
	.A(FE_RN_271_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_316_0 (
	.Y(FE_RN_270_0),
	.A(a[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_315_0 (
	.Y(FE_RN_269_0),
	.A(\u_div/SumTmp[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X4M FE_RC_314_0 (
	.Y(\u_div/PartRem[4][1] ),
	.S0(quotient[4]),
	.B(FE_RN_269_0),
	.A(FE_RN_270_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_313_0 (
	.Y(FE_RN_268_0),
	.A(a[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_312_0 (
	.Y(FE_RN_267_0),
	.B(n18),
	.A(FE_RN_268_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B1X8M FE_RC_311_0 (
	.Y(FE_RN_266_0),
	.B0(FE_RN_267_0),
	.A1N(a[4]),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X8M FE_RC_310_0 (
	.Y(FE_RN_265_0),
	.B(\u_div/CryTmp[3][1] ),
	.A(FE_RN_266_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_309_0 (
	.Y(FE_RN_264_0),
	.A(FE_RN_250_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X6M FE_RC_308_0 (
	.Y(FE_RN_263_0),
	.B(FE_RN_264_0),
	.A(FE_RN_253_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_307_0 (
	.Y(FE_RN_262_0),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX4M FE_RC_306_0 (
	.Y(FE_RN_261_0),
	.B(FE_RN_262_0),
	.AN(\u_div/CryTmp[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX8M FE_RC_305_0 (
	.Y(FE_RN_260_0),
	.B(FE_RN_261_0),
	.AN(FE_RN_253_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_304_0 (
	.Y(FE_RN_259_0),
	.A(\u_div/SumTmp[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X6M FE_RC_303_0 (
	.Y(FE_RN_258_0),
	.S0(FE_RN_259_0),
	.B(FE_RN_260_0),
	.A(FE_RN_263_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_302_0 (
	.Y(FE_RN_257_0),
	.B(quotient[4]),
	.A(FE_RN_258_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B1X4M FE_RC_301_0 (
	.Y(\u_div/SumTmp[3][1] ),
	.B0(FE_RN_257_0),
	.A1N(FE_RN_265_0),
	.A0(quotient[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_300_0 (
	.Y(FE_RN_256_0),
	.A(a[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX8M FE_RC_299_0 (
	.Y(FE_RN_255_0),
	.B(FE_RN_256_0),
	.AN(FE_RN_250_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_298_0 (
	.Y(FE_RN_254_0),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX8M FE_RC_297_0 (
	.Y(FE_RN_253_0),
	.B(FE_RN_254_0),
	.AN(\u_div/CryTmp[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_296_0 (
	.Y(FE_RN_252_0),
	.A(FE_RN_253_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_295_0 (
	.Y(FE_RN_251_0),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX8M FE_RC_294_0 (
	.Y(FE_RN_250_0),
	.B(FE_RN_251_0),
	.AN(\u_div/CryTmp[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_293_0 (
	.Y(FE_RN_249_0),
	.A(\u_div/SumTmp[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX8M FE_RC_292_0 (
	.Y(FE_RN_248_0),
	.B(FE_RN_249_0),
	.AN(FE_RN_250_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_291_0 (
	.Y(FE_RN_247_0),
	.B(quotient[4]),
	.A(FE_RN_248_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B11X4M FE_RC_290_0 (
	.Y(\u_div/CryTmp[3][2] ),
	.C0(FE_RN_247_0),
	.B0(FE_RN_252_0),
	.A1N(FE_RN_255_0),
	.A0(quotient[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_243_0 (
	.Y(FE_RN_205_0),
	.A(\u_div/CryTmp[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X2M FE_RC_242_0 (
	.Y(FE_RN_204_0),
	.B(n16),
	.A(\u_div/PartRem[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_241_0 (
	.Y(FE_RN_203_0),
	.B(n16),
	.A(\u_div/PartRem[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_240_0 (
	.Y(FE_RN_202_0),
	.B(FE_RN_198_0),
	.A(FE_RN_203_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_239_0 (
	.Y(FE_RN_201_0),
	.B(\u_div/CryTmp[4][3] ),
	.A(FE_RN_202_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M FE_RC_238_0 (
	.Y(\u_div/SumTmp[4][3] ),
	.B0(FE_RN_201_0),
	.A1N(FE_RN_204_0),
	.A0N(FE_RN_205_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X1M FE_RC_237_0 (
	.Y(FE_RN_200_0),
	.C(n21),
	.B(n16),
	.A(\u_div/PartRem[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_236_0 (
	.Y(FE_RN_199_0),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX4M FE_RC_235_0 (
	.Y(FE_RN_198_0),
	.B(FE_RN_199_0),
	.AN(\u_div/PartRem[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M FE_RC_234_0 (
	.Y(FE_RN_197_0),
	.C(n21),
	.B(\u_div/CryTmp[4][3] ),
	.A(FE_RN_198_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_201_0 (
	.Y(FE_RN_168_0),
	.B(\u_div/PartRem[6][1] ),
	.A(FE_RN_155_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X5M FE_RC_200_0 (
	.Y(\u_div/CryTmp[5][2] ),
	.B(FE_RN_168_0),
	.A(FE_RN_157_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X3M FE_RC_199_0 (
	.Y(FE_RN_167_0),
	.B(FE_RN_161_0),
	.A(FE_RN_151_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X5M FE_RC_198_0 (
	.Y(quotient[5]),
	.B(FE_RN_119_0),
	.A(FE_RN_167_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M FE_RC_197_0 (
	.Y(FE_RN_166_0),
	.B1(\u_div/CryTmp[5][1] ),
	.B0(n18),
	.A1N(n18),
	.A0N(\u_div/CryTmp[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M FE_RC_196_0 (
	.Y(FE_RN_165_0),
	.B0(\u_div/PartRem[6][1] ),
	.A1N(FE_RN_155_0),
	.A0N(FE_RN_157_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M FE_RC_195_0 (
	.Y(\u_div/SumTmp[5][1] ),
	.B0(FE_RN_165_0),
	.A1(\u_div/PartRem[6][1] ),
	.A0(FE_RN_166_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_194_0 (
	.Y(FE_RN_164_0),
	.A(FE_RN_98_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_193_0 (
	.Y(FE_RN_163_0),
	.B(FE_RN_164_0),
	.A(FE_RN_161_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_192_0 (
	.Y(FE_RN_162_0),
	.A(FE_RN_157_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X4M FE_RC_191_0 (
	.Y(FE_RN_161_0),
	.B1(FE_RN_162_0),
	.B0(n20),
	.A1N(FE_RN_154_0),
	.A0(\u_div/PartRem[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_190_0 (
	.Y(FE_RN_160_0),
	.B(FE_RN_105_0),
	.A(FE_RN_161_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X3M FE_RC_189_0 (
	.Y(FE_RN_159_0),
	.C(FE_RN_119_0),
	.B(FE_RN_163_0),
	.A(FE_RN_160_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X3M FE_RC_188_0 (
	.Y(FE_RN_158_0),
	.B(\u_div/SumTmp[5][0] ),
	.A(FE_RN_159_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_187_0 (
	.Y(FE_RN_157_0),
	.B(\u_div/CryTmp[5][1] ),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_186_0 (
	.Y(FE_RN_156_0),
	.A(FE_RN_157_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M FE_RC_185_0 (
	.Y(FE_RN_155_0),
	.B(\u_div/CryTmp[5][1] ),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_184_0 (
	.Y(FE_RN_154_0),
	.B(n20),
	.A(FE_RN_155_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X4M FE_RC_183_0 (
	.Y(FE_RN_153_0),
	.B0(FE_RN_154_0),
	.A1N(\u_div/PartRem[6][1] ),
	.A0N(FE_RN_156_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_182_0 (
	.Y(FE_RN_152_0),
	.A(FE_RN_105_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X3M FE_RC_181_0 (
	.Y(FE_RN_151_0),
	.B(FE_RN_98_0),
	.A(FE_RN_152_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_180_0 (
	.Y(FE_RN_150_0),
	.B(FE_RN_153_0),
	.A(FE_RN_151_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M FE_RC_179_0 (
	.Y(FE_RN_149_0),
	.C(FE_RN_119_0),
	.B(a[5]),
	.A(FE_RN_150_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X5M FE_RC_178_0 (
	.Y(\u_div/PartRem[5][1] ),
	.B(FE_RN_158_0),
	.A(FE_RN_149_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX4M FE_RC_177_0 (
	.Y(FE_RN_39_0),
	.C(FE_RN_40_0),
	.B(FE_RN_36_0),
	.AN(FE_RN_43_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX3M FE_RC_176_0 (
	.Y(quotient[6]),
	.A(FE_RN_100_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_175_0 (
	.Y(FE_RN_148_0),
	.A(FE_RN_118_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_174_0 (
	.Y(FE_RN_147_0),
	.A(FE_RN_100_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_173_0 (
	.Y(FE_RN_146_0),
	.A(FE_RN_7_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_172_0 (
	.Y(FE_RN_145_0),
	.A(FE_RN_104_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_171_0 (
	.Y(FE_RN_144_0),
	.A(FE_RN_115_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_170_0 (
	.Y(FE_RN_143_0),
	.A(FE_RN_7_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X4M FE_RC_169_0 (
	.Y(FE_RN_142_0),
	.B0(FE_RN_109_0),
	.A1(FE_RN_143_0),
	.A0(FE_RN_144_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M FE_RC_168_0 (
	.Y(FE_RN_141_0),
	.B0(FE_RN_142_0),
	.A1N(FE_RN_145_0),
	.A0N(FE_RN_146_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X3M FE_RC_167_0 (
	.Y(FE_RN_140_0),
	.B(FE_RN_147_0),
	.A(FE_RN_141_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_166_0 (
	.Y(\u_div/PartRem[6][2] ),
	.B(FE_RN_148_0),
	.A(FE_RN_140_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_165_0 (
	.Y(FE_RN_139_0),
	.A(FE_RN_100_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X4M FE_RC_164_0 (
	.Y(FE_RN_138_0),
	.C(\u_div/PartRem[7][1] ),
	.B(FE_RN_128_0),
	.A(FE_RN_139_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X4M FE_RC_163_0 (
	.Y(FE_RN_137_0),
	.B0(FE_RN_138_0),
	.A1(FE_RN_128_0),
	.A0(FE_RN_112_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_162_0 (
	.Y(FE_RN_136_0),
	.A(FE_RN_100_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_161_0 (
	.Y(FE_RN_135_0),
	.A(FE_RN_104_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X5M FE_RC_160_0 (
	.Y(FE_RN_134_0),
	.B(FE_RN_128_0),
	.A(FE_RN_122_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X4M FE_RC_159_0 (
	.Y(FE_RN_133_0),
	.B0(FE_RN_134_0),
	.A1(FE_RN_128_0),
	.A0(FE_RN_135_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_158_0 (
	.Y(FE_RN_132_0),
	.A(FE_RN_20_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_157_0 (
	.Y(FE_RN_131_0),
	.A(FE_RN_20_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_156_0 (
	.Y(FE_RN_130_0),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_155_0 (
	.Y(FE_RN_129_0),
	.B(\u_div/CryTmp[5][2] ),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B1X8M FE_RC_154_0 (
	.Y(FE_RN_128_0),
	.B0(FE_RN_129_0),
	.A1N(FE_RN_130_0),
	.A0(\u_div/CryTmp[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X4M FE_RC_153_0 (
	.Y(FE_RN_127_0),
	.B(FE_RN_131_0),
	.A(FE_RN_128_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X4M FE_RC_152_0 (
	.Y(FE_RN_126_0),
	.B0(FE_RN_127_0),
	.A1(FE_RN_132_0),
	.A0(FE_RN_128_0), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X2M FE_RC_151_0 (
	.Y(FE_RN_125_0),
	.S0(FE_RN_7_0),
	.B(FE_RN_126_0),
	.A(FE_RN_133_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X3M FE_RC_150_0 (
	.Y(FE_RN_124_0),
	.B(FE_RN_136_0),
	.A(FE_RN_125_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_149_0 (
	.Y(\u_div/SumTmp[5][2] ),
	.B(FE_RN_137_0),
	.A(FE_RN_124_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_148_0 (
	.Y(FE_RN_123_0),
	.A(FE_RN_118_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_147_0 (
	.Y(FE_RN_122_0),
	.B(FE_RN_115_0),
	.A(FE_RN_104_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_146_0 (
	.Y(FE_RN_121_0),
	.B(FE_RN_122_0),
	.A(FE_RN_99_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B11X4M FE_RC_145_0 (
	.Y(FE_RN_120_0),
	.C0(FE_RN_121_0),
	.B0(FE_RN_123_0),
	.A1N(FE_RN_109_0),
	.A0(FE_RN_100_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M FE_RC_144_0 (
	.Y(FE_RN_119_0),
	.C(n20),
	.B(n17),
	.A(FE_RN_120_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKAND2X8M FE_RC_143_0 (
	.Y(FE_RN_118_0),
	.B(\u_div/PartRem[7][1] ),
	.A(FE_RN_100_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_142_0 (
	.Y(FE_RN_117_0),
	.A(FE_RN_118_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_141_0 (
	.Y(FE_RN_116_0),
	.A(FE_RN_28_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX4M FE_RC_140_0 (
	.Y(FE_RN_115_0),
	.B(FE_RN_26_0),
	.AN(FE_RN_116_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_139_0 (
	.Y(FE_RN_114_0),
	.A(FE_RN_115_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_138_0 (
	.Y(FE_RN_113_0),
	.B(FE_RN_114_0),
	.A(FE_RN_99_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_137_0 (
	.Y(FE_RN_112_0),
	.B(FE_RN_117_0),
	.A(FE_RN_113_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_136_0 (
	.Y(FE_RN_111_0),
	.A(FE_RN_112_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_135_0 (
	.Y(FE_RN_110_0),
	.A(FE_RN_7_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X4M FE_RC_134_0 (
	.Y(FE_RN_109_0),
	.B(FE_RN_110_0),
	.A(FE_RN_20_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_133_0 (
	.Y(FE_RN_108_0),
	.A(FE_RN_109_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X6M FE_RC_132_0 (
	.Y(FE_RN_107_0),
	.B(FE_RN_100_0),
	.A(FE_RN_108_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X4M FE_RC_131_0 (
	.Y(FE_RN_106_0),
	.B(n17),
	.A(FE_RN_107_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_130_0 (
	.Y(FE_RN_105_0),
	.B(FE_RN_111_0),
	.A(FE_RN_106_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_129_0 (
	.Y(FE_RN_104_0),
	.B(FE_RN_11_0),
	.A(FE_RN_29_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_128_0 (
	.Y(FE_RN_103_0),
	.A(FE_RN_104_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_127_0 (
	.Y(FE_RN_102_0),
	.A(FE_RN_45_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX4M FE_RC_126_0 (
	.Y(FE_RN_101_0),
	.C(FE_RN_40_0),
	.B(FE_RN_36_0),
	.AN(FE_RN_43_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X6M FE_RC_125_0 (
	.Y(FE_RN_100_0),
	.B(FE_RN_102_0),
	.A(FE_RN_101_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X8M FE_RC_124_0 (
	.Y(FE_RN_99_0),
	.B(FE_RN_7_0),
	.A(FE_RN_100_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_123_0 (
	.Y(FE_RN_98_0),
	.B(FE_RN_103_0),
	.A(FE_RN_99_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X6M FE_RC_70_0 (
	.Y(FE_RN_7_0),
	.D(FE_RN_9_0),
	.C(n21),
	.B(\u_div/CryTmp[7][1] ),
	.A(FE_RN_8_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_68_0 (
	.Y(FE_RN_51_0),
	.A(FE_RN_45_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_67_0 (
	.Y(FE_RN_50_0),
	.A(FE_RN_10_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M FE_RC_66_0 (
	.Y(FE_RN_49_0),
	.C(FE_RN_13_0),
	.B(FE_RN_50_0),
	.A(FE_RN_41_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M FE_RC_65_0 (
	.Y(FE_RN_48_0),
	.C(FE_RN_17_0),
	.B(FE_RN_36_0),
	.A(FE_RN_49_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_64_0 (
	.Y(FE_RN_47_0),
	.B(FE_RN_51_0),
	.A(FE_RN_48_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_63_0 (
	.Y(FE_RN_46_0),
	.B(a[6]),
	.A(FE_RN_47_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X5M FE_RC_62_0 (
	.Y(FE_RN_45_0),
	.B(n17),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_61_0 (
	.Y(FE_RN_44_0),
	.A(FE_RN_45_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_60_0 (
	.Y(FE_RN_43_0),
	.A(FE_RN_17_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_59_0 (
	.Y(FE_RN_42_0),
	.A(FE_RN_10_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X4M FE_RC_58_0 (
	.Y(FE_RN_41_0),
	.D(FE_RN_8_0),
	.C(FE_RN_9_0),
	.B(\u_div/CryTmp[7][1] ),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M FE_RC_57_0 (
	.Y(FE_RN_40_0),
	.C(FE_RN_13_0),
	.B(FE_RN_42_0),
	.A(FE_RN_41_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M FE_RC_55_0 (
	.Y(FE_RN_38_0),
	.C(\u_div/SumTmp[6][0] ),
	.B(FE_RN_44_0),
	.A(FE_RN_39_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_54_0 (
	.Y(\u_div/PartRem[6][1] ),
	.B(FE_RN_46_0),
	.A(FE_RN_38_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X4M FE_RC_52_0 (
	.Y(FE_RN_37_0),
	.D(FE_RN_9_0),
	.C(n21),
	.B(\u_div/CryTmp[7][1] ),
	.A(FE_RN_8_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M FE_RC_51_0 (
	.Y(FE_RN_36_0),
	.C(FE_RN_37_0),
	.B(FE_RN_13_0),
	.A(FE_RN_15_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_48_0 (
	.Y(FE_RN_34_0),
	.A(FE_RN_11_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_47_0 (
	.Y(FE_RN_33_0),
	.A(FE_RN_10_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_46_0 (
	.Y(FE_RN_32_0),
	.B(FE_RN_7_0),
	.A(FE_RN_33_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B1X4M FE_RC_45_0 (
	.Y(\u_div/PartRem[7][1] ),
	.B0(FE_RN_32_0),
	.A1N(FE_RN_34_0),
	.A0(FE_RN_7_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_44_0 (
	.Y(FE_RN_31_0),
	.A(FE_RN_18_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M FE_RC_43_0 (
	.Y(FE_RN_30_0),
	.B0(FE_RN_31_0),
	.A1(\u_div/CryTmp[6][1] ),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_42_0 (
	.Y(FE_RN_29_0),
	.A(FE_RN_30_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_41_0 (
	.Y(FE_RN_28_0),
	.A(FE_RN_11_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_40_0 (
	.Y(FE_RN_27_0),
	.A(FE_RN_18_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X3M FE_RC_39_0 (
	.Y(FE_RN_26_0),
	.B(FE_RN_13_0),
	.A(FE_RN_27_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_37_0 (
	.Y(FE_RN_24_0),
	.A(\u_div/CryTmp[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_36_0 (
	.Y(FE_RN_23_0),
	.A(\u_div/CryTmp[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X8M FE_RC_35_0 (
	.Y(FE_RN_22_0),
	.B1(n18),
	.B0(FE_RN_10_0),
	.A1N(FE_RN_10_0),
	.A0N(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X3M FE_RC_34_0 (
	.Y(FE_RN_21_0),
	.B(FE_RN_23_0),
	.A(FE_RN_22_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X4M FE_RC_33_0 (
	.Y(FE_RN_20_0),
	.B0(FE_RN_21_0),
	.A1(FE_RN_24_0),
	.A0(FE_RN_22_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_31_0 (
	.Y(FE_RN_19_0),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX8M FE_RC_30_0 (
	.Y(FE_RN_18_0),
	.B(FE_RN_19_0),
	.AN(\u_div/CryTmp[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_29_0 (
	.Y(FE_RN_17_0),
	.A(FE_RN_18_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_27_0 (
	.Y(FE_RN_15_0),
	.A(FE_RN_11_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_26_0 (
	.Y(FE_RN_14_0),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX8M FE_RC_25_0 (
	.Y(FE_RN_13_0),
	.B(FE_RN_14_0),
	.AN(\u_div/CryTmp[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M FE_RC_22_0 (
	.Y(quotient[7]),
	.A(FE_RN_7_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_21_0 (
	.Y(FE_RN_11_0),
	.A(\u_div/SumTmp[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_20_0 (
	.Y(FE_RN_10_0),
	.A(a[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_19_0 (
	.Y(FE_RN_9_0),
	.A(FE_RN_4_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X4M FE_RC_18_0 (
	.Y(FE_RN_8_0),
	.B(FE_RN_5_0),
	.A(FE_RN_1_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X6M FE_RC_15_0 (
	.Y(n21),
	.C(FE_RN_0_0),
	.B(n15),
	.A(FE_RN_2_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_14_0 (
	.Y(FE_RN_6_0),
	.A(FE_RN_1_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X8M FE_RC_13_0 (
	.Y(n20),
	.B(FE_RN_6_0),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_12_0 (
	.Y(FE_RN_5_0),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_11_0 (
	.Y(FE_RN_4_0),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X12M FE_RC_8_0 (
	.Y(n22),
	.B(b[7]),
	.A(b[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X8M FE_RC_7_0 (
	.Y(FE_RN_2_0),
	.B(b[7]),
	.A(b[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX8M FE_RC_5_0 (
	.Y(FE_RN_1_0),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX10M FE_RC_3_0 (
	.Y(n14),
	.A(b[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_2_0 (
	.Y(FE_RN_0_0),
	.A(b[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX10M FE_RC_0_0 (
	.Y(n15),
	.A(b[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX2M \u_div/u_fa_PartRem_0_0_5  (
	.CO(\u_div/CryTmp[0][6] ),
	.CI(\u_div/CryTmp[0][5] ),
	.B(n14),
	.A(\u_div/PartRem[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX2M \u_div/u_fa_PartRem_0_0_6  (
	.CO(\u_div/CryTmp[0][7] ),
	.CI(\u_div/CryTmp[0][6] ),
	.B(n163),
	.A(\u_div/PartRem[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX2M \u_div/u_fa_PartRem_0_0_7  (
	.CO(quotient[0]),
	.CI(\u_div/CryTmp[0][7] ),
	.B(n12),
	.A(\u_div/PartRem[1][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX1M \u_div/u_fa_PartRem_0_0_1  (
	.CO(\u_div/CryTmp[0][2] ),
	.CI(\u_div/CryTmp[0][1] ),
	.B(n18),
	.A(\u_div/PartRem[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX1M \u_div/u_fa_PartRem_0_4_1  (
	.S(\u_div/SumTmp[4][1] ),
	.CO(\u_div/CryTmp[4][2] ),
	.CI(\u_div/CryTmp[4][1] ),
	.B(n18),
	.A(\u_div/PartRem[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX2M \u_div/u_fa_PartRem_0_0_2  (
	.CO(\u_div/CryTmp[0][3] ),
	.CI(\u_div/CryTmp[0][2] ),
	.B(n17),
	.A(\u_div/PartRem[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX2M \u_div/u_fa_PartRem_0_0_3  (
	.CO(\u_div/CryTmp[0][4] ),
	.CI(\u_div/CryTmp[0][3] ),
	.B(n16),
	.A(\u_div/PartRem[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX2M \u_div/u_fa_PartRem_0_0_4  (
	.CO(\u_div/CryTmp[0][5] ),
	.CI(\u_div/CryTmp[0][4] ),
	.B(n15),
	.A(\u_div/PartRem[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX1M \u_div/u_fa_PartRem_0_4_2  (
	.S(\u_div/SumTmp[4][2] ),
	.CO(\u_div/CryTmp[4][3] ),
	.CI(\u_div/CryTmp[4][2] ),
	.B(n17),
	.A(\u_div/PartRem[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX12M U1 (
	.Y(n19),
	.A(b[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U2 (
	.Y(\u_div/SumTmp[7][0] ),
	.B(a[7]),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U3 (
	.Y(\u_div/SumTmp[6][0] ),
	.B(a[6]),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U4 (
	.Y(\u_div/SumTmp[5][0] ),
	.B(a[5]),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U5 (
	.Y(\u_div/SumTmp[4][0] ),
	.B(a[4]),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U6 (
	.Y(\u_div/SumTmp[3][0] ),
	.B(a[3]),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U7 (
	.Y(\u_div/SumTmp[2][0] ),
	.B(a[2]),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U8 (
	.Y(\u_div/CryTmp[7][1] ),
	.B(a[7]),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U9 (
	.Y(\u_div/SumTmp[1][0] ),
	.B(a[1]),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX12M U10 (
	.Y(n18),
	.A(b[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X1M U11 (
	.Y(\u_div/CryTmp[5][1] ),
	.B(n3),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U12 (
	.Y(n3),
	.A(a[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U13 (
	.Y(n2),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U14 (
	.Y(\u_div/CryTmp[4][1] ),
	.B(n5),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U15 (
	.Y(n5),
	.A(a[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U16 (
	.Y(n4),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U17 (
	.Y(\u_div/CryTmp[3][1] ),
	.B(n7),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U18 (
	.Y(n7),
	.A(a[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U19 (
	.Y(n6),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U20 (
	.Y(\u_div/CryTmp[2][1] ),
	.B(n9),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U21 (
	.Y(n9),
	.A(a[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U22 (
	.Y(n8),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U23 (
	.Y(\u_div/CryTmp[1][1] ),
	.B(n183),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U25 (
	.Y(\u_div/CryTmp[0][1] ),
	.B(n184),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U27 (
	.Y(\u_div/CryTmp[6][1] ),
	.B(n1),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U28 (
	.Y(n1),
	.A(a[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX12M U30 (
	.Y(n17),
	.A(b[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX6M U31 (
	.Y(n16),
	.A(b[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U34 (
	.Y(n12),
	.A(b[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U35 (
	.Y(\u_div/PartRem[1][7] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][6] ),
	.A(\u_div/PartRem[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U36 (
	.Y(\u_div/PartRem[2][6] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][5] ),
	.A(\u_div/PartRem[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U37 (
	.Y(\u_div/PartRem[3][5] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][4] ),
	.A(\u_div/PartRem[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U38 (
	.Y(\u_div/PartRem[4][4] ),
	.S0(quotient[4]),
	.B(\u_div/SumTmp[4][3] ),
	.A(\u_div/PartRem[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X6M U39 (
	.Y(\u_div/PartRem[5][3] ),
	.S0(quotient[5]),
	.B(\u_div/SumTmp[5][2] ),
	.A(\u_div/PartRem[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U42 (
	.Y(\u_div/PartRem[1][6] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][5] ),
	.A(\u_div/PartRem[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U43 (
	.Y(\u_div/PartRem[2][5] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][4] ),
	.A(\u_div/PartRem[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U44 (
	.Y(\u_div/PartRem[3][4] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][3] ),
	.A(\u_div/PartRem[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U46 (
	.Y(\u_div/PartRem[5][2] ),
	.S0(quotient[5]),
	.B(\u_div/SumTmp[5][1] ),
	.A(\u_div/PartRem[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U48 (
	.Y(\u_div/PartRem[1][5] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][4] ),
	.A(\u_div/PartRem[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U49 (
	.Y(\u_div/PartRem[2][4] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][3] ),
	.A(\u_div/PartRem[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X8M U50 (
	.Y(\u_div/PartRem[3][3] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][2] ),
	.A(\u_div/PartRem[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U53 (
	.Y(\u_div/PartRem[1][4] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][3] ),
	.A(\u_div/PartRem[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U54 (
	.Y(\u_div/PartRem[2][3] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][2] ),
	.A(\u_div/PartRem[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U57 (
	.Y(\u_div/PartRem[1][3] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][2] ),
	.A(\u_div/PartRem[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U60 (
	.Y(\u_div/PartRem[1][2] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][1] ),
	.A(\u_div/PartRem[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module bit16_alu_DW01_sub_0 (
	A, 
	B, 
	CI, 
	DIFF, 
	CO, 
	n160, 
	n161, 
	n162, 
	n186, 
	n185, 
	n184, 
	n187, 
	n163, 
	VDD, 
	VSS);
   input [8:0] A;
   input [8:0] B;
   input CI;
   output [8:0] DIFF;
   output CO;
   input n160;
   input n161;
   input n162;
   input n186;
   input n185;
   input n184;
   input n187;
   input n163;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n2;
   wire [9:0] carry;

   // Module instantiations
   ADDFX2M U2_7 (
	.S(DIFF[7]),
	.CO(carry[8]),
	.CI(carry[7]),
	.B(n2),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_5 (
	.S(DIFF[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(n185),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_4 (
	.S(DIFF[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(n186),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_3 (
	.S(DIFF[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(n162),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_2 (
	.S(DIFF[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(n161),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_1 (
	.S(DIFF[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(n187),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_6 (
	.S(DIFF[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(n163),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U1 (
	.Y(DIFF[0]),
	.B(A[0]),
	.A(n160), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U4 (
	.Y(carry[1]),
	.B(n184),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U11 (
	.Y(n2),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U12 (
	.Y(DIFF[8]),
	.A(carry[8]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module bit16_alu_DW01_add_0 (
	A, 
	B, 
	CI, 
	SUM, 
	CO, 
	VDD, 
	VSS);
   input [8:0] A;
   input [8:0] B;
   input CI;
   output [8:0] SUM;
   output CO;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire [8:1] carry;

   // Module instantiations
   ADDFX2M U1_7 (
	.S(SUM[7]),
	.CO(SUM[8]),
	.CI(carry[7]),
	.B(B[7]),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.CI(n1),
	.B(B[1]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(B[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(B[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(B[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(B[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(B[6]),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U1 (
	.Y(n1),
	.B(A[0]),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U2 (
	.Y(SUM[0]),
	.B(A[0]),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module bit16_alu_DW02_mult_0 (
	A, 
	B, 
	TC, 
	PRODUCT, 
	n160, 
	n161, 
	n162, 
	n184, 
	n183, 
	n182, 
	n181, 
	n180, 
	n179, 
	n178, 
	n177, 
	n187, 
	n163, 
	n185, 
	n186, 
	VDD, 
	VSS);
   input [7:0] A;
   input [7:0] B;
   input TC;
   output [15:0] PRODUCT;
   input n160;
   input n161;
   input n162;
   input n184;
   input n183;
   input n182;
   input n181;
   input n180;
   input n179;
   input n178;
   input n177;
   input n187;
   input n163;
   input n185;
   input n186;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \ab[7][7] ;
   wire \ab[7][6] ;
   wire \ab[7][5] ;
   wire \ab[7][4] ;
   wire \ab[7][3] ;
   wire \ab[7][2] ;
   wire \ab[7][1] ;
   wire \ab[7][0] ;
   wire \ab[6][7] ;
   wire \ab[6][6] ;
   wire \ab[6][5] ;
   wire \ab[6][4] ;
   wire \ab[6][3] ;
   wire \ab[6][2] ;
   wire \ab[6][1] ;
   wire \ab[6][0] ;
   wire \ab[5][7] ;
   wire \ab[5][6] ;
   wire \ab[5][5] ;
   wire \ab[5][4] ;
   wire \ab[5][3] ;
   wire \ab[5][2] ;
   wire \ab[5][1] ;
   wire \ab[5][0] ;
   wire \ab[4][7] ;
   wire \ab[4][6] ;
   wire \ab[4][5] ;
   wire \ab[4][4] ;
   wire \ab[4][3] ;
   wire \ab[4][2] ;
   wire \ab[4][1] ;
   wire \ab[4][0] ;
   wire \ab[3][7] ;
   wire \ab[3][6] ;
   wire \ab[3][5] ;
   wire \ab[3][4] ;
   wire \ab[3][3] ;
   wire \ab[3][2] ;
   wire \ab[3][1] ;
   wire \ab[3][0] ;
   wire \ab[2][7] ;
   wire \ab[2][6] ;
   wire \ab[2][5] ;
   wire \ab[2][4] ;
   wire \ab[2][3] ;
   wire \ab[2][2] ;
   wire \ab[2][1] ;
   wire \ab[2][0] ;
   wire \ab[1][7] ;
   wire \ab[1][6] ;
   wire \ab[1][5] ;
   wire \ab[1][4] ;
   wire \ab[1][3] ;
   wire \ab[1][2] ;
   wire \ab[1][1] ;
   wire \ab[1][0] ;
   wire \ab[0][7] ;
   wire \ab[0][6] ;
   wire \ab[0][5] ;
   wire \ab[0][4] ;
   wire \ab[0][3] ;
   wire \ab[0][2] ;
   wire \ab[0][1] ;
   wire \CARRYB[7][6] ;
   wire \CARRYB[7][5] ;
   wire \CARRYB[7][4] ;
   wire \CARRYB[7][3] ;
   wire \CARRYB[7][2] ;
   wire \CARRYB[7][1] ;
   wire \CARRYB[7][0] ;
   wire \CARRYB[6][6] ;
   wire \CARRYB[6][5] ;
   wire \CARRYB[6][4] ;
   wire \CARRYB[6][3] ;
   wire \CARRYB[6][2] ;
   wire \CARRYB[6][1] ;
   wire \CARRYB[6][0] ;
   wire \CARRYB[5][6] ;
   wire \CARRYB[5][5] ;
   wire \CARRYB[5][4] ;
   wire \CARRYB[5][3] ;
   wire \CARRYB[5][2] ;
   wire \CARRYB[5][1] ;
   wire \CARRYB[5][0] ;
   wire \CARRYB[4][6] ;
   wire \CARRYB[4][5] ;
   wire \CARRYB[4][4] ;
   wire \CARRYB[4][3] ;
   wire \CARRYB[4][2] ;
   wire \CARRYB[4][1] ;
   wire \CARRYB[4][0] ;
   wire \CARRYB[3][6] ;
   wire \CARRYB[3][5] ;
   wire \CARRYB[3][4] ;
   wire \CARRYB[3][3] ;
   wire \CARRYB[3][2] ;
   wire \CARRYB[3][1] ;
   wire \CARRYB[3][0] ;
   wire \CARRYB[2][6] ;
   wire \CARRYB[2][5] ;
   wire \CARRYB[2][4] ;
   wire \CARRYB[2][3] ;
   wire \CARRYB[2][2] ;
   wire \CARRYB[2][1] ;
   wire \CARRYB[2][0] ;
   wire \SUMB[7][6] ;
   wire \SUMB[7][5] ;
   wire \SUMB[7][4] ;
   wire \SUMB[7][3] ;
   wire \SUMB[7][2] ;
   wire \SUMB[7][1] ;
   wire \SUMB[7][0] ;
   wire \SUMB[6][6] ;
   wire \SUMB[6][5] ;
   wire \SUMB[6][4] ;
   wire \SUMB[6][3] ;
   wire \SUMB[6][2] ;
   wire \SUMB[6][1] ;
   wire \SUMB[5][6] ;
   wire \SUMB[5][5] ;
   wire \SUMB[5][4] ;
   wire \SUMB[5][3] ;
   wire \SUMB[5][2] ;
   wire \SUMB[5][1] ;
   wire \SUMB[4][6] ;
   wire \SUMB[4][5] ;
   wire \SUMB[4][4] ;
   wire \SUMB[4][3] ;
   wire \SUMB[4][2] ;
   wire \SUMB[4][1] ;
   wire \SUMB[3][6] ;
   wire \SUMB[3][5] ;
   wire \SUMB[3][4] ;
   wire \SUMB[3][3] ;
   wire \SUMB[3][2] ;
   wire \SUMB[3][1] ;
   wire \SUMB[2][6] ;
   wire \SUMB[2][5] ;
   wire \SUMB[2][4] ;
   wire \SUMB[2][3] ;
   wire \SUMB[2][2] ;
   wire \SUMB[2][1] ;
   wire \SUMB[1][6] ;
   wire \SUMB[1][5] ;
   wire \SUMB[1][4] ;
   wire \SUMB[1][3] ;
   wire \SUMB[1][2] ;
   wire \SUMB[1][1] ;
   wire \A1[12] ;
   wire \A1[11] ;
   wire \A1[10] ;
   wire \A1[9] ;
   wire \A1[8] ;
   wire \A1[7] ;
   wire \A1[6] ;
   wire \A1[4] ;
   wire \A1[3] ;
   wire \A1[2] ;
   wire \A1[1] ;
   wire \A1[0] ;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n33;

   // Module instantiations
   ADDFX2M S1_6_0 (
	.S(\A1[4] ),
	.CO(\CARRYB[6][0] ),
	.CI(\SUMB[5][1] ),
	.B(\CARRYB[5][0] ),
	.A(\ab[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_4 (
	.S(\SUMB[6][4] ),
	.CO(\CARRYB[6][4] ),
	.CI(\SUMB[5][5] ),
	.B(\CARRYB[5][4] ),
	.A(\ab[6][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_3 (
	.S(\SUMB[6][3] ),
	.CO(\CARRYB[6][3] ),
	.CI(\SUMB[5][4] ),
	.B(\CARRYB[5][3] ),
	.A(\ab[6][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_2 (
	.S(\SUMB[6][2] ),
	.CO(\CARRYB[6][2] ),
	.CI(\SUMB[5][3] ),
	.B(\CARRYB[5][2] ),
	.A(\ab[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_5_0 (
	.S(\A1[3] ),
	.CO(\CARRYB[5][0] ),
	.CI(\SUMB[4][1] ),
	.B(\CARRYB[4][0] ),
	.A(\ab[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_5 (
	.S(\SUMB[6][5] ),
	.CO(\CARRYB[6][5] ),
	.CI(\SUMB[5][6] ),
	.B(\CARRYB[5][5] ),
	.A(\ab[6][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_4 (
	.S(\SUMB[5][4] ),
	.CO(\CARRYB[5][4] ),
	.CI(\SUMB[4][5] ),
	.B(\CARRYB[4][4] ),
	.A(\ab[5][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_3 (
	.S(\SUMB[5][3] ),
	.CO(\CARRYB[5][3] ),
	.CI(\SUMB[4][4] ),
	.B(\CARRYB[4][3] ),
	.A(\ab[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_2 (
	.S(\SUMB[5][2] ),
	.CO(\CARRYB[5][2] ),
	.CI(\SUMB[4][3] ),
	.B(\CARRYB[4][2] ),
	.A(\ab[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_4_0 (
	.S(\A1[2] ),
	.CO(\CARRYB[4][0] ),
	.CI(\SUMB[3][1] ),
	.B(\CARRYB[3][0] ),
	.A(\ab[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_5 (
	.S(\SUMB[5][5] ),
	.CO(\CARRYB[5][5] ),
	.CI(\SUMB[4][6] ),
	.B(\CARRYB[4][5] ),
	.A(\ab[5][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_4 (
	.S(\SUMB[4][4] ),
	.CO(\CARRYB[4][4] ),
	.CI(\SUMB[3][5] ),
	.B(\CARRYB[3][4] ),
	.A(\ab[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_3 (
	.S(\SUMB[4][3] ),
	.CO(\CARRYB[4][3] ),
	.CI(\SUMB[3][4] ),
	.B(\CARRYB[3][3] ),
	.A(\ab[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_2 (
	.S(\SUMB[4][2] ),
	.CO(\CARRYB[4][2] ),
	.CI(\SUMB[3][3] ),
	.B(\CARRYB[3][2] ),
	.A(\ab[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_3_0 (
	.S(\A1[1] ),
	.CO(\CARRYB[3][0] ),
	.CI(\SUMB[2][1] ),
	.B(\CARRYB[2][0] ),
	.A(\ab[3][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_5 (
	.S(\SUMB[4][5] ),
	.CO(\CARRYB[4][5] ),
	.CI(\SUMB[3][6] ),
	.B(\CARRYB[3][5] ),
	.A(\ab[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_4 (
	.S(\SUMB[3][4] ),
	.CO(\CARRYB[3][4] ),
	.CI(\SUMB[2][5] ),
	.B(\CARRYB[2][4] ),
	.A(\ab[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_3 (
	.S(\SUMB[3][3] ),
	.CO(\CARRYB[3][3] ),
	.CI(\SUMB[2][4] ),
	.B(\CARRYB[2][3] ),
	.A(\ab[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_2 (
	.S(\SUMB[3][2] ),
	.CO(\CARRYB[3][2] ),
	.CI(\SUMB[2][3] ),
	.B(\CARRYB[2][2] ),
	.A(\ab[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_5 (
	.S(\SUMB[3][5] ),
	.CO(\CARRYB[3][5] ),
	.CI(\SUMB[2][6] ),
	.B(\CARRYB[2][5] ),
	.A(\ab[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_6_6 (
	.S(\SUMB[6][6] ),
	.CO(\CARRYB[6][6] ),
	.CI(\ab[5][7] ),
	.B(\CARRYB[5][6] ),
	.A(\ab[6][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_5_6 (
	.S(\SUMB[5][6] ),
	.CO(\CARRYB[5][6] ),
	.CI(\ab[4][7] ),
	.B(\CARRYB[4][6] ),
	.A(\ab[5][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_4_6 (
	.S(\SUMB[4][6] ),
	.CO(\CARRYB[4][6] ),
	.CI(\ab[3][7] ),
	.B(\CARRYB[3][6] ),
	.A(\ab[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_3_6 (
	.S(\SUMB[3][6] ),
	.CO(\CARRYB[3][6] ),
	.CI(\ab[2][7] ),
	.B(\CARRYB[2][6] ),
	.A(\ab[3][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_2_6 (
	.S(\SUMB[2][6] ),
	.CO(\CARRYB[2][6] ),
	.CI(\ab[1][7] ),
	.B(n9),
	.A(\ab[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_2_0 (
	.S(\A1[0] ),
	.CO(\CARRYB[2][0] ),
	.CI(\SUMB[1][1] ),
	.B(n8),
	.A(\ab[2][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_4 (
	.S(\SUMB[2][4] ),
	.CO(\CARRYB[2][4] ),
	.CI(\SUMB[1][5] ),
	.B(n7),
	.A(\ab[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_3 (
	.S(\SUMB[2][3] ),
	.CO(\CARRYB[2][3] ),
	.CI(\SUMB[1][4] ),
	.B(n6),
	.A(\ab[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_2 (
	.S(\SUMB[2][2] ),
	.CO(\CARRYB[2][2] ),
	.CI(\SUMB[1][3] ),
	.B(n5),
	.A(\ab[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_5 (
	.S(\SUMB[2][5] ),
	.CO(\CARRYB[2][5] ),
	.CI(\SUMB[1][6] ),
	.B(n4),
	.A(\ab[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_0 (
	.S(\SUMB[7][0] ),
	.CO(\CARRYB[7][0] ),
	.CI(\SUMB[6][1] ),
	.B(\CARRYB[6][0] ),
	.A(\ab[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S5_6 (
	.S(\SUMB[7][6] ),
	.CO(\CARRYB[7][6] ),
	.CI(\ab[6][7] ),
	.B(\CARRYB[6][6] ),
	.A(\ab[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_4 (
	.S(\SUMB[7][4] ),
	.CO(\CARRYB[7][4] ),
	.CI(\SUMB[6][5] ),
	.B(\CARRYB[6][4] ),
	.A(\ab[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_3 (
	.S(\SUMB[7][3] ),
	.CO(\CARRYB[7][3] ),
	.CI(\SUMB[6][4] ),
	.B(\CARRYB[6][3] ),
	.A(\ab[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_2 (
	.S(\SUMB[7][2] ),
	.CO(\CARRYB[7][2] ),
	.CI(\SUMB[6][3] ),
	.B(\CARRYB[6][2] ),
	.A(\ab[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_5 (
	.S(\SUMB[7][5] ),
	.CO(\CARRYB[7][5] ),
	.CI(\SUMB[6][6] ),
	.B(\CARRYB[6][5] ),
	.A(\ab[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_1 (
	.S(\SUMB[6][1] ),
	.CO(\CARRYB[6][1] ),
	.CI(\SUMB[5][2] ),
	.B(\CARRYB[5][1] ),
	.A(\ab[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_1 (
	.S(\SUMB[5][1] ),
	.CO(\CARRYB[5][1] ),
	.CI(\SUMB[4][2] ),
	.B(\CARRYB[4][1] ),
	.A(\ab[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_1 (
	.S(\SUMB[4][1] ),
	.CO(\CARRYB[4][1] ),
	.CI(\SUMB[3][2] ),
	.B(\CARRYB[3][1] ),
	.A(\ab[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_1 (
	.S(\SUMB[3][1] ),
	.CO(\CARRYB[3][1] ),
	.CI(\SUMB[2][2] ),
	.B(\CARRYB[2][1] ),
	.A(\ab[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_1 (
	.S(\SUMB[2][1] ),
	.CO(\CARRYB[2][1] ),
	.CI(\SUMB[1][2] ),
	.B(n3),
	.A(\ab[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_1 (
	.S(\SUMB[7][1] ),
	.CO(\CARRYB[7][1] ),
	.CI(\SUMB[6][2] ),
	.B(\CARRYB[6][1] ),
	.A(\ab[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U2 (
	.Y(n3),
	.B(\ab[1][1] ),
	.A(\ab[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U3 (
	.Y(n4),
	.B(\ab[1][5] ),
	.A(\ab[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U4 (
	.Y(n5),
	.B(\ab[1][2] ),
	.A(\ab[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U5 (
	.Y(n6),
	.B(\ab[1][3] ),
	.A(\ab[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U6 (
	.Y(n7),
	.B(\ab[1][4] ),
	.A(\ab[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U7 (
	.Y(n8),
	.B(\ab[1][0] ),
	.A(\ab[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U8 (
	.Y(n9),
	.B(\ab[1][6] ),
	.A(\ab[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U9 (
	.Y(n10),
	.B(\ab[7][7] ),
	.A(\CARRYB[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U10 (
	.Y(n23),
	.A(\ab[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U11 (
	.Y(\A1[7] ),
	.B(\SUMB[7][2] ),
	.A(\CARRYB[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U12 (
	.Y(\A1[12] ),
	.B(\ab[7][7] ),
	.A(\CARRYB[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U13 (
	.Y(\A1[8] ),
	.B(\SUMB[7][3] ),
	.A(\CARRYB[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U14 (
	.Y(\A1[10] ),
	.B(\SUMB[7][5] ),
	.A(\CARRYB[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U15 (
	.Y(\A1[9] ),
	.B(\SUMB[7][4] ),
	.A(\CARRYB[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U16 (
	.Y(\A1[11] ),
	.B(\SUMB[7][6] ),
	.A(\CARRYB[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U17 (
	.Y(n24),
	.A(\ab[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U18 (
	.Y(n21),
	.A(\ab[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U19 (
	.Y(n22),
	.A(\ab[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n20),
	.A(\ab[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U21 (
	.Y(n19),
	.A(\ab[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U22 (
	.Y(\SUMB[1][2] ),
	.B(n20),
	.A(\ab[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U23 (
	.Y(\A1[6] ),
	.B(n17),
	.A(\CARRYB[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U24 (
	.Y(n17),
	.A(\SUMB[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U25 (
	.Y(n11),
	.B(\SUMB[7][1] ),
	.A(\CARRYB[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U26 (
	.Y(n12),
	.B(\SUMB[7][2] ),
	.A(\CARRYB[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U27 (
	.Y(n13),
	.B(\SUMB[7][4] ),
	.A(\CARRYB[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U28 (
	.Y(n14),
	.B(\SUMB[7][6] ),
	.A(\CARRYB[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U29 (
	.Y(n15),
	.B(\SUMB[7][3] ),
	.A(\CARRYB[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U30 (
	.Y(n16),
	.B(\SUMB[7][5] ),
	.A(\CARRYB[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U31 (
	.Y(\SUMB[1][6] ),
	.B(n24),
	.A(\ab[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U32 (
	.Y(\SUMB[1][3] ),
	.B(n21),
	.A(\ab[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U33 (
	.Y(\SUMB[1][4] ),
	.B(n22),
	.A(\ab[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U34 (
	.Y(\SUMB[1][5] ),
	.B(n23),
	.A(\ab[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U35 (
	.Y(\SUMB[1][1] ),
	.B(n19),
	.A(\ab[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U46 (
	.Y(PRODUCT[1]),
	.B(n18),
	.A(\ab[1][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U47 (
	.Y(n18),
	.A(\ab[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U53 (
	.Y(n33),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U55 (
	.Y(\ab[7][7] ),
	.B(n33),
	.A(n177), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U56 (
	.Y(\ab[7][6] ),
	.B(n163),
	.A(n177), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U57 (
	.Y(\ab[7][5] ),
	.B(n185),
	.A(n177), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U58 (
	.Y(\ab[7][4] ),
	.B(n186),
	.A(n177), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U59 (
	.Y(\ab[7][3] ),
	.B(n162),
	.A(n177), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U60 (
	.Y(\ab[7][2] ),
	.B(n161),
	.A(n177), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U61 (
	.Y(\ab[7][1] ),
	.B(n187),
	.A(n177), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U62 (
	.Y(\ab[7][0] ),
	.B(n160),
	.A(n177), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U63 (
	.Y(\ab[6][7] ),
	.B(n178),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U64 (
	.Y(\ab[6][6] ),
	.B(n178),
	.A(n163), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U65 (
	.Y(\ab[6][5] ),
	.B(n178),
	.A(n185), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U66 (
	.Y(\ab[6][4] ),
	.B(n178),
	.A(n186), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U67 (
	.Y(\ab[6][3] ),
	.B(n178),
	.A(n162), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U68 (
	.Y(\ab[6][2] ),
	.B(n178),
	.A(n161), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U69 (
	.Y(\ab[6][1] ),
	.B(n178),
	.A(n187), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U70 (
	.Y(\ab[6][0] ),
	.B(n178),
	.A(n160), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U71 (
	.Y(\ab[5][7] ),
	.B(n179),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U72 (
	.Y(\ab[5][6] ),
	.B(n179),
	.A(n163), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U73 (
	.Y(\ab[5][5] ),
	.B(n179),
	.A(n185), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U74 (
	.Y(\ab[5][4] ),
	.B(n179),
	.A(n186), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U75 (
	.Y(\ab[5][3] ),
	.B(n179),
	.A(n162), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U76 (
	.Y(\ab[5][2] ),
	.B(n179),
	.A(n161), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U77 (
	.Y(\ab[5][1] ),
	.B(n179),
	.A(n187), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U78 (
	.Y(\ab[5][0] ),
	.B(n179),
	.A(n160), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U79 (
	.Y(\ab[4][7] ),
	.B(n180),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U80 (
	.Y(\ab[4][6] ),
	.B(n180),
	.A(n163), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U81 (
	.Y(\ab[4][5] ),
	.B(n180),
	.A(n185), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U82 (
	.Y(\ab[4][4] ),
	.B(n180),
	.A(n186), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U83 (
	.Y(\ab[4][3] ),
	.B(n180),
	.A(n162), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U84 (
	.Y(\ab[4][2] ),
	.B(n180),
	.A(n161), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U85 (
	.Y(\ab[4][1] ),
	.B(n180),
	.A(n187), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U86 (
	.Y(\ab[4][0] ),
	.B(n180),
	.A(n160), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U87 (
	.Y(\ab[3][7] ),
	.B(n181),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U88 (
	.Y(\ab[3][6] ),
	.B(n181),
	.A(n163), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U89 (
	.Y(\ab[3][5] ),
	.B(n181),
	.A(n185), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U90 (
	.Y(\ab[3][4] ),
	.B(n181),
	.A(n186), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U91 (
	.Y(\ab[3][3] ),
	.B(n181),
	.A(n162), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U92 (
	.Y(\ab[3][2] ),
	.B(n181),
	.A(n161), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U93 (
	.Y(\ab[3][1] ),
	.B(n181),
	.A(n187), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U94 (
	.Y(\ab[3][0] ),
	.B(n181),
	.A(n160), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U95 (
	.Y(\ab[2][7] ),
	.B(n182),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U96 (
	.Y(\ab[2][6] ),
	.B(n182),
	.A(n163), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U97 (
	.Y(\ab[2][5] ),
	.B(n182),
	.A(n185), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U98 (
	.Y(\ab[2][4] ),
	.B(n182),
	.A(n186), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U99 (
	.Y(\ab[2][3] ),
	.B(n182),
	.A(n162), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U100 (
	.Y(\ab[2][2] ),
	.B(n182),
	.A(n161), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U101 (
	.Y(\ab[2][1] ),
	.B(n182),
	.A(n187), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U102 (
	.Y(\ab[2][0] ),
	.B(n182),
	.A(n160), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U103 (
	.Y(\ab[1][7] ),
	.B(n183),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U104 (
	.Y(\ab[1][6] ),
	.B(n183),
	.A(n163), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U105 (
	.Y(\ab[1][5] ),
	.B(n183),
	.A(n185), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U106 (
	.Y(\ab[1][4] ),
	.B(n183),
	.A(n186), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U107 (
	.Y(\ab[1][3] ),
	.B(n183),
	.A(n162), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U108 (
	.Y(\ab[1][2] ),
	.B(n183),
	.A(n161), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U109 (
	.Y(\ab[1][1] ),
	.B(n183),
	.A(n187), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U110 (
	.Y(\ab[1][0] ),
	.B(n183),
	.A(n160), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U111 (
	.Y(\ab[0][7] ),
	.B(n184),
	.A(n33), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U112 (
	.Y(\ab[0][6] ),
	.B(n184),
	.A(n163), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U113 (
	.Y(\ab[0][5] ),
	.B(n184),
	.A(n185), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U114 (
	.Y(\ab[0][4] ),
	.B(n184),
	.A(n186), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U115 (
	.Y(\ab[0][3] ),
	.B(n184),
	.A(n162), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U116 (
	.Y(\ab[0][2] ),
	.B(n184),
	.A(n161), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U117 (
	.Y(\ab[0][1] ),
	.B(n184),
	.A(n187), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U118 (
	.Y(PRODUCT[0]),
	.B(n184),
	.A(n160), 
	.VDD(VDD), 
	.VSS(VSS));
   bit16_alu_DW01_add_1 FS_1 (
	.A({ 1'b0,
		\A1[12] ,
		\A1[11] ,
		\A1[10] ,
		\A1[9] ,
		\A1[8] ,
		\A1[7] ,
		\A1[6] ,
		\SUMB[7][0] ,
		\A1[4] ,
		\A1[3] ,
		\A1[2] ,
		\A1[1] ,
		\A1[0]  }),
	.B({ n10,
		n14,
		n16,
		n13,
		n15,
		n12,
		n11,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0 }),
	.CI(1'b0),
	.SUM({ PRODUCT[15],
		PRODUCT[14],
		PRODUCT[13],
		PRODUCT[12],
		PRODUCT[11],
		PRODUCT[10],
		PRODUCT[9],
		PRODUCT[8],
		PRODUCT[7],
		PRODUCT[6],
		PRODUCT[5],
		PRODUCT[4],
		PRODUCT[3],
		PRODUCT[2] }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module bit16_alu_DW01_add_1 (
	A, 
	B, 
	CI, 
	SUM, 
	CO, 
	VDD, 
	VSS);
   input [13:0] A;
   input [13:0] B;
   input CI;
   output [13:0] SUM;
   output CO;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;

   // Module instantiations
   NAND2X2M U2 (
	.Y(n15),
	.B(B[7]),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21BX2M U3 (
	.Y(n1),
	.B0N(n19),
	.A1(A[12]),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U4 (
	.Y(n9),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U5 (
	.Y(SUM[7]),
	.B(n8),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U6 (
	.Y(n8),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U7 (
	.Y(SUM[13]),
	.B(n1),
	.A(B[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U8 (
	.Y(SUM[6]),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U9 (
	.Y(SUM[0]),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U10 (
	.Y(SUM[1]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U11 (
	.Y(SUM[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U12 (
	.Y(SUM[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U13 (
	.Y(SUM[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U14 (
	.Y(SUM[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U15 (
	.Y(SUM[9]),
	.B(n11),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U16 (
	.Y(n11),
	.B(n13),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U17 (
	.Y(SUM[8]),
	.B(n15),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U18 (
	.Y(n14),
	.B(n17),
	.AN(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U19 (
	.Y(n19),
	.B0(B[12]),
	.A1(n18),
	.A0(A[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U20 (
	.Y(SUM[12]),
	.C(n18),
	.B(A[12]),
	.A(B[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21BX1M U21 (
	.Y(n18),
	.B0N(n22),
	.A1(n21),
	.A0(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U22 (
	.Y(SUM[11]),
	.B(n23),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U23 (
	.Y(n23),
	.B(n20),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U24 (
	.Y(n20),
	.B(A[11]),
	.A(B[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U25 (
	.Y(n22),
	.B(A[11]),
	.A(B[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X1M U26 (
	.Y(n21),
	.B0(n26),
	.A1(n25),
	.A0(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U27 (
	.Y(SUM[10]),
	.B(n25),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X1M U28 (
	.Y(n25),
	.B0(n12),
	.A1N(n13),
	.A0N(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U29 (
	.Y(n12),
	.B(A[9]),
	.A(B[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U30 (
	.Y(n13),
	.B(A[9]),
	.A(B[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X1M U31 (
	.Y(n10),
	.B0(n17),
	.A1(n16),
	.A0(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U32 (
	.Y(n17),
	.B(A[8]),
	.A(B[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U33 (
	.Y(n16),
	.B(A[8]),
	.A(B[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U34 (
	.Y(n27),
	.B(n26),
	.AN(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U35 (
	.Y(n26),
	.B(A[10]),
	.A(B[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U36 (
	.Y(n24),
	.B(A[10]),
	.A(B[10]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module fifo_top_test_1 (
	w_clk, 
	w_rst_n, 
	rd_clk, 
	rd_rst_n, 
	w_inc, 
	rd_inc, 
	w_data, 
	rd_data, 
	full_flag, 
	empty_flag, 
	test_si3, 
	test_si2, 
	test_si1, 
	test_so3, 
	test_so2, 
	test_so1, 
	test_se, 
	FE_OFN3_scan_rst_sync1_mux_out, 
	FE_OFN4_scan_rst_sync1_mux_out, 
	scan_clk_ref_clk_mux_out__L4_N1, 
	VDD, 
	VSS);
   input w_clk;
   input w_rst_n;
   input rd_clk;
   input rd_rst_n;
   input w_inc;
   input rd_inc;
   input [7:0] w_data;
   output [7:0] rd_data;
   output full_flag;
   output empty_flag;
   input test_si3;
   input test_si2;
   input test_si1;
   output test_so3;
   output test_so2;
   output test_so1;
   input test_se;
   input FE_OFN3_scan_rst_sync1_mux_out;
   input FE_OFN4_scan_rst_sync1_mux_out;
   input scan_clk_ref_clk_mux_out__L4_N1;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_UNCONNECTED_0;
   wire n5;
   wire n6;
   wire n9;
   wire [4:0] sync_grey_coded_rd_ptr;
   wire [4:0] wr_ptr_grey_coded;
   wire [3:0] w_address;
   wire [3:0] rd_address;
   wire [4:0] sync_grey_coded_wr_ptr;
   wire [4:0] rd_ptr_grey_coded;

   assign test_so3 = sync_grey_coded_wr_ptr[4] ;

   // Module instantiations
   full_gen_test_1 dut1 (
	.sync_grey_coded_rd_ptr({ sync_grey_coded_rd_ptr[4],
		sync_grey_coded_rd_ptr[3],
		sync_grey_coded_rd_ptr[2],
		sync_grey_coded_rd_ptr[1],
		sync_grey_coded_rd_ptr[0] }),
	.w_clk(scan_clk_ref_clk_mux_out__L4_N1),
	.w_rst_n(w_rst_n),
	.w_inc(w_inc),
	.wr_ptr_grey_coded({ wr_ptr_grey_coded[4],
		wr_ptr_grey_coded[3],
		wr_ptr_grey_coded[2],
		wr_ptr_grey_coded[1],
		wr_ptr_grey_coded[0] }),
	.w_address({ w_address[3],
		w_address[2],
		w_address[1],
		w_address[0] }),
	.full_flag(full_flag),
	.test_si(test_si1),
	.test_so(n9),
	.test_se(test_se),
	.FE_OFN4_scan_rst_sync1_mux_out(FE_OFN4_scan_rst_sync1_mux_out), 
	.VDD(VDD), 
	.VSS(VSS));
   fifo_memory_test_1 dut2 (
	.w_clk(scan_clk_ref_clk_mux_out__L4_N1),
	.w_rst_n(w_rst_n),
	.rd_clk(rd_clk),
	.rd_rst_n(FE_UNCONNECTED_0),
	.w_address({ w_address[3],
		w_address[2],
		w_address[1],
		w_address[0] }),
	.rd_address({ rd_address[3],
		rd_address[2],
		rd_address[1],
		rd_address[0] }),
	.w_inc(w_inc),
	.full_flag(full_flag),
	.w_data({ w_data[7],
		w_data[6],
		w_data[5],
		w_data[4],
		w_data[3],
		w_data[2],
		w_data[1],
		w_data[0] }),
	.rd_data({ rd_data[7],
		rd_data[6],
		rd_data[5],
		rd_data[4],
		rd_data[3],
		rd_data[2],
		rd_data[1],
		rd_data[0] }),
	.test_si3(test_si3),
	.test_si2(test_si2),
	.test_si1(n9),
	.test_so3(n6),
	.test_so2(test_so2),
	.test_so1(test_so1),
	.test_se(test_se),
	.FE_OFN3_scan_rst_sync1_mux_out(FE_OFN3_scan_rst_sync1_mux_out),
	.FE_OFN4_scan_rst_sync1_mux_out(FE_OFN4_scan_rst_sync1_mux_out), 
	.VDD(VDD), 
	.VSS(VSS));
   empty_gen_test_1 dut3 (
	.sync_grey_coded_wr_ptr({ sync_grey_coded_wr_ptr[4],
		sync_grey_coded_wr_ptr[3],
		sync_grey_coded_wr_ptr[2],
		sync_grey_coded_wr_ptr[1],
		sync_grey_coded_wr_ptr[0] }),
	.rd_clk(rd_clk),
	.rd_rst_n(rd_rst_n),
	.rd_inc(rd_inc),
	.rd_ptr_grey_coded({ rd_ptr_grey_coded[4],
		rd_ptr_grey_coded[3],
		rd_ptr_grey_coded[2],
		rd_ptr_grey_coded[1],
		rd_ptr_grey_coded[0] }),
	.rd_address({ rd_address[3],
		rd_address[2],
		rd_address[1],
		rd_address[0] }),
	.empty_flag(empty_flag),
	.test_si(n6),
	.test_so(n5),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   synchronizer_test_0 dut4 (
	.d1({ rd_ptr_grey_coded[4],
		rd_ptr_grey_coded[3],
		rd_ptr_grey_coded[2],
		rd_ptr_grey_coded[1],
		rd_ptr_grey_coded[0] }),
	.clk(w_clk),
	.rst_n(w_rst_n),
	.q2({ sync_grey_coded_rd_ptr[4],
		sync_grey_coded_rd_ptr[3],
		sync_grey_coded_rd_ptr[2],
		sync_grey_coded_rd_ptr[1],
		sync_grey_coded_rd_ptr[0] }),
	.test_si(n5),
	.test_se(test_se),
	.scan_clk_ref_clk_mux_out__L4_N1(scan_clk_ref_clk_mux_out__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   synchronizer_test_1 dut5 (
	.d1({ wr_ptr_grey_coded[4],
		wr_ptr_grey_coded[3],
		wr_ptr_grey_coded[2],
		wr_ptr_grey_coded[1],
		wr_ptr_grey_coded[0] }),
	.clk(rd_clk),
	.rst_n(rd_rst_n),
	.q2({ sync_grey_coded_wr_ptr[4],
		sync_grey_coded_wr_ptr[3],
		sync_grey_coded_wr_ptr[2],
		sync_grey_coded_wr_ptr[1],
		sync_grey_coded_wr_ptr[0] }),
	.test_si(sync_grey_coded_rd_ptr[4]),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module full_gen_test_1 (
	sync_grey_coded_rd_ptr, 
	w_clk, 
	w_rst_n, 
	w_inc, 
	wr_ptr_grey_coded, 
	w_address, 
	full_flag, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN4_scan_rst_sync1_mux_out, 
	VDD, 
	VSS);
   input [4:0] sync_grey_coded_rd_ptr;
   input w_clk;
   input w_rst_n;
   input w_inc;
   output [4:0] wr_ptr_grey_coded;
   output [3:0] w_address;
   output full_flag;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN4_scan_rst_sync1_mux_out;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N11;
   wire N12;
   wire N13;
   wire N14;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire \add_21/carry[4] ;
   wire \add_21/carry[3] ;
   wire \add_21/carry[2] ;
   wire n10;
   wire [4:0] wr_ptr;

   assign test_so = wr_ptr[4] ;

   // Module instantiations
   SDFFRQX2M \w_address_reg[3]  (
	.SI(w_address[2]),
	.SE(test_se),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(w_address[3]),
	.D(n25),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \w_address_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(w_rst_n),
	.Q(w_address[0]),
	.D(n28),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \w_address_reg[2]  (
	.SI(w_address[1]),
	.SE(test_se),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(w_address[2]),
	.D(n26),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \w_address_reg[1]  (
	.SI(w_address[0]),
	.SE(test_se),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(w_address[1]),
	.D(n27),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \wr_ptr_reg[4]  (
	.SI(wr_ptr[3]),
	.SE(test_se),
	.RN(w_rst_n),
	.Q(wr_ptr[4]),
	.D(n29),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \wr_ptr_reg[0]  (
	.SI(w_address[3]),
	.SE(test_se),
	.RN(w_rst_n),
	.Q(wr_ptr[0]),
	.D(n30),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \wr_ptr_reg[3]  (
	.SI(wr_ptr[2]),
	.SE(test_se),
	.RN(w_rst_n),
	.Q(wr_ptr[3]),
	.D(n22),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \wr_ptr_reg[2]  (
	.SI(wr_ptr[1]),
	.SE(test_se),
	.RN(w_rst_n),
	.Q(wr_ptr[2]),
	.D(n23),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \wr_ptr_reg[1]  (
	.SI(wr_ptr[0]),
	.SE(test_se),
	.RN(w_rst_n),
	.Q(wr_ptr[1]),
	.D(n24),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U12 (
	.Y(n10),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U13 (
	.Y(n11),
	.B(n15),
	.A(w_inc), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U14 (
	.Y(full_flag),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U15 (
	.Y(n26),
	.B(n13),
	.A(w_address[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U16 (
	.Y(n15),
	.D(n19),
	.C(n18),
	.B(n17),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U17 (
	.Y(n16),
	.B(sync_grey_coded_rd_ptr[0]),
	.A(wr_ptr_grey_coded[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U18 (
	.Y(n17),
	.B(sync_grey_coded_rd_ptr[1]),
	.A(wr_ptr_grey_coded[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U19 (
	.Y(n19),
	.B(sync_grey_coded_rd_ptr[2]),
	.A(wr_ptr_grey_coded[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U20 (
	.Y(n13),
	.B(n14),
	.A(w_address[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U21 (
	.Y(n18),
	.B(n21),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U22 (
	.Y(n20),
	.B(sync_grey_coded_rd_ptr[4]),
	.A(wr_ptr_grey_coded[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U23 (
	.Y(n21),
	.B(sync_grey_coded_rd_ptr[3]),
	.A(wr_ptr_grey_coded[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U24 (
	.Y(n14),
	.B(n10),
	.A(w_address[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U25 (
	.Y(n24),
	.B1(n11),
	.B0(wr_ptr[1]),
	.A1(n10),
	.A0(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U26 (
	.Y(n23),
	.B1(n11),
	.B0(wr_ptr[2]),
	.A1(n10),
	.A0(N12), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U27 (
	.Y(n22),
	.B1(n11),
	.B0(wr_ptr[3]),
	.A1(n10),
	.A0(N13), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U28 (
	.Y(n29),
	.B1(n11),
	.B0(wr_ptr[4]),
	.A1(n10),
	.A0(N14), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U29 (
	.Y(n30),
	.B1(n11),
	.B0(wr_ptr[0]),
	.A1N(wr_ptr[0]),
	.A0(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U30 (
	.Y(n25),
	.B(n12),
	.A(w_address[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U31 (
	.Y(n12),
	.B(n13),
	.AN(w_address[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U32 (
	.Y(n27),
	.B(n14),
	.A(w_address[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U33 (
	.Y(n28),
	.B(n10),
	.A(w_address[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U34 (
	.S(N11),
	.CO(\add_21/carry[2] ),
	.B(wr_ptr[0]),
	.A(wr_ptr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U35 (
	.S(N12),
	.CO(\add_21/carry[3] ),
	.B(\add_21/carry[2] ),
	.A(wr_ptr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U36 (
	.S(N13),
	.CO(\add_21/carry[4] ),
	.B(\add_21/carry[3] ),
	.A(wr_ptr[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U37 (
	.Y(N14),
	.B(wr_ptr[4]),
	.A(\add_21/carry[4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   grey_code_gen_0 wr_ptr_gc (
	.binary_data({ wr_ptr[4],
		wr_ptr[3],
		wr_ptr[2],
		wr_ptr[1],
		wr_ptr[0] }),
	.grey_coded_data({ wr_ptr_grey_coded[4],
		wr_ptr_grey_coded[3],
		wr_ptr_grey_coded[2],
		wr_ptr_grey_coded[1],
		wr_ptr_grey_coded[0] }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module grey_code_gen_0 (
	binary_data, 
	grey_coded_data, 
	VDD, 
	VSS);
   input [4:0] binary_data;
   output [4:0] grey_coded_data;
   inout VDD;
   inout VSS;

   // Module instantiations
   CLKXOR2X2M U1 (
	.Y(grey_coded_data[0]),
	.B(binary_data[0]),
	.A(binary_data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U2 (
	.Y(grey_coded_data[1]),
	.B(binary_data[1]),
	.A(binary_data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U3 (
	.Y(grey_coded_data[2]),
	.B(binary_data[2]),
	.A(binary_data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U4 (
	.Y(grey_coded_data[3]),
	.B(binary_data[3]),
	.A(binary_data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U5 (
	.Y(grey_coded_data[4]),
	.A(binary_data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module fifo_memory_test_1 (
	w_clk, 
	w_rst_n, 
	rd_clk, 
	rd_rst_n, 
	w_address, 
	rd_address, 
	w_inc, 
	full_flag, 
	w_data, 
	rd_data, 
	test_si3, 
	test_si2, 
	test_si1, 
	test_so3, 
	test_so2, 
	test_so1, 
	test_se, 
	FE_OFN3_scan_rst_sync1_mux_out, 
	FE_OFN4_scan_rst_sync1_mux_out, 
	VDD, 
	VSS);
   input w_clk;
   input w_rst_n;
   input rd_clk;
   input rd_rst_n;
   input [3:0] w_address;
   input [3:0] rd_address;
   input w_inc;
   input full_flag;
   input [7:0] w_data;
   output [7:0] rd_data;
   input test_si3;
   input test_si2;
   input test_si1;
   output test_so3;
   output test_so2;
   output test_so1;
   input test_se;
   input FE_OFN3_scan_rst_sync1_mux_out;
   input FE_OFN4_scan_rst_sync1_mux_out;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_OFN9_SO_4_;
   wire FE_OFN8_SO_3_;
   wire N9;
   wire N10;
   wire N11;
   wire N12;
   wire \fifo[0][7] ;
   wire \fifo[0][6] ;
   wire \fifo[0][5] ;
   wire \fifo[0][4] ;
   wire \fifo[0][3] ;
   wire \fifo[0][2] ;
   wire \fifo[0][1] ;
   wire \fifo[0][0] ;
   wire \fifo[1][7] ;
   wire \fifo[1][6] ;
   wire \fifo[1][5] ;
   wire \fifo[1][4] ;
   wire \fifo[1][3] ;
   wire \fifo[1][2] ;
   wire \fifo[1][1] ;
   wire \fifo[1][0] ;
   wire \fifo[2][7] ;
   wire \fifo[2][6] ;
   wire \fifo[2][5] ;
   wire \fifo[2][4] ;
   wire \fifo[2][3] ;
   wire \fifo[2][2] ;
   wire \fifo[2][1] ;
   wire \fifo[2][0] ;
   wire \fifo[3][7] ;
   wire \fifo[3][6] ;
   wire \fifo[3][5] ;
   wire \fifo[3][4] ;
   wire \fifo[3][3] ;
   wire \fifo[3][2] ;
   wire \fifo[3][1] ;
   wire \fifo[3][0] ;
   wire \fifo[4][7] ;
   wire \fifo[4][6] ;
   wire \fifo[4][5] ;
   wire \fifo[4][4] ;
   wire \fifo[4][3] ;
   wire \fifo[4][2] ;
   wire \fifo[4][1] ;
   wire \fifo[4][0] ;
   wire \fifo[5][7] ;
   wire \fifo[5][6] ;
   wire \fifo[5][5] ;
   wire \fifo[5][4] ;
   wire \fifo[5][3] ;
   wire \fifo[5][2] ;
   wire \fifo[5][1] ;
   wire \fifo[5][0] ;
   wire \fifo[6][7] ;
   wire \fifo[6][6] ;
   wire \fifo[6][5] ;
   wire \fifo[6][4] ;
   wire \fifo[6][3] ;
   wire \fifo[6][2] ;
   wire \fifo[6][1] ;
   wire \fifo[6][0] ;
   wire \fifo[7][7] ;
   wire \fifo[7][6] ;
   wire \fifo[7][5] ;
   wire \fifo[7][4] ;
   wire \fifo[7][3] ;
   wire \fifo[7][2] ;
   wire \fifo[7][1] ;
   wire \fifo[7][0] ;
   wire \fifo[8][7] ;
   wire \fifo[8][6] ;
   wire \fifo[8][5] ;
   wire \fifo[8][4] ;
   wire \fifo[8][3] ;
   wire \fifo[8][2] ;
   wire \fifo[8][1] ;
   wire \fifo[8][0] ;
   wire \fifo[9][7] ;
   wire \fifo[9][6] ;
   wire \fifo[9][5] ;
   wire \fifo[9][4] ;
   wire \fifo[9][3] ;
   wire \fifo[9][2] ;
   wire \fifo[9][1] ;
   wire \fifo[9][0] ;
   wire \fifo[10][7] ;
   wire \fifo[10][6] ;
   wire \fifo[10][5] ;
   wire \fifo[10][4] ;
   wire \fifo[10][3] ;
   wire \fifo[10][2] ;
   wire \fifo[10][1] ;
   wire \fifo[10][0] ;
   wire \fifo[11][7] ;
   wire \fifo[11][6] ;
   wire \fifo[11][5] ;
   wire \fifo[11][4] ;
   wire \fifo[11][3] ;
   wire \fifo[11][2] ;
   wire \fifo[11][1] ;
   wire \fifo[11][0] ;
   wire \fifo[12][7] ;
   wire \fifo[12][6] ;
   wire \fifo[12][5] ;
   wire \fifo[12][4] ;
   wire \fifo[12][3] ;
   wire \fifo[12][2] ;
   wire \fifo[12][1] ;
   wire \fifo[12][0] ;
   wire \fifo[13][7] ;
   wire \fifo[13][6] ;
   wire \fifo[13][5] ;
   wire \fifo[13][4] ;
   wire \fifo[13][3] ;
   wire \fifo[13][2] ;
   wire \fifo[13][1] ;
   wire \fifo[13][0] ;
   wire \fifo[14][7] ;
   wire \fifo[14][6] ;
   wire \fifo[14][5] ;
   wire \fifo[14][4] ;
   wire \fifo[14][3] ;
   wire \fifo[14][2] ;
   wire \fifo[14][1] ;
   wire \fifo[14][0] ;
   wire \fifo[15][7] ;
   wire \fifo[15][6] ;
   wire \fifo[15][5] ;
   wire \fifo[15][4] ;
   wire \fifo[15][3] ;
   wire \fifo[15][2] ;
   wire \fifo[15][1] ;
   wire \fifo[15][0] ;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n318;
   wire n319;
   wire n321;
   wire n322;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;

   assign N9 = rd_address[0] ;
   assign N10 = rd_address[1] ;
   assign N11 = rd_address[2] ;
   assign N12 = rd_address[3] ;
   assign test_so1 = \fifo[5][0]  ;
   assign test_so3 = \fifo[15][7]  ;
   assign test_so2 = \fifo[15][2]  ;

   // Module instantiations
   BUFX10M FE_OFC9_SO_4_ (
	.Y(\fifo[5][0] ),
	.A(FE_OFN9_SO_4_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX10M FE_OFC8_SO_3_ (
	.Y(\fifo[15][2] ),
	.A(FE_OFN8_SO_3_), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[1][7]  (
	.SI(\fifo[1][6] ),
	.SE(n355),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[1][7] ),
	.D(n286),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[1][6]  (
	.SI(\fifo[1][5] ),
	.SE(n358),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[1][6] ),
	.D(n285),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[1][5]  (
	.SI(\fifo[1][4] ),
	.SE(n357),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[1][5] ),
	.D(n284),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[1][4]  (
	.SI(\fifo[1][3] ),
	.SE(n356),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[1][4] ),
	.D(n283),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[1][3]  (
	.SI(\fifo[1][2] ),
	.SE(n355),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[1][3] ),
	.D(n282),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[1][2]  (
	.SI(\fifo[1][1] ),
	.SE(n358),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[1][2] ),
	.D(n281),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[1][1]  (
	.SI(\fifo[1][0] ),
	.SE(n357),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[1][1] ),
	.D(n280),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[1][0]  (
	.SI(\fifo[0][7] ),
	.SE(n356),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[1][0] ),
	.D(n279),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[5][7]  (
	.SI(\fifo[5][6] ),
	.SE(n355),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[5][7] ),
	.D(n254),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[5][6]  (
	.SI(\fifo[5][5] ),
	.SE(n358),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[5][6] ),
	.D(n253),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[5][5]  (
	.SI(\fifo[5][4] ),
	.SE(n357),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[5][5] ),
	.D(n252),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[5][4]  (
	.SI(\fifo[5][3] ),
	.SE(n356),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[5][4] ),
	.D(n251),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[5][3]  (
	.SI(\fifo[5][2] ),
	.SE(n355),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[5][3] ),
	.D(n250),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[5][2]  (
	.SI(\fifo[5][1] ),
	.SE(n358),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[5][2] ),
	.D(n249),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[5][1]  (
	.SI(test_si2),
	.SE(n357),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[5][1] ),
	.D(n248),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[9][7]  (
	.SI(\fifo[9][6] ),
	.SE(n355),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[9][7] ),
	.D(n222),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[9][6]  (
	.SI(\fifo[9][5] ),
	.SE(n358),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[9][6] ),
	.D(n221),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[9][5]  (
	.SI(\fifo[9][4] ),
	.SE(n357),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[9][5] ),
	.D(n220),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[9][4]  (
	.SI(\fifo[9][3] ),
	.SE(n356),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[9][4] ),
	.D(n219),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[9][3]  (
	.SI(\fifo[9][2] ),
	.SE(n355),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[9][3] ),
	.D(n218),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[9][2]  (
	.SI(\fifo[9][1] ),
	.SE(n358),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[9][2] ),
	.D(n217),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[9][1]  (
	.SI(\fifo[9][0] ),
	.SE(n357),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[9][1] ),
	.D(n216),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[9][0]  (
	.SI(\fifo[8][7] ),
	.SE(n356),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[9][0] ),
	.D(n215),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[13][7]  (
	.SI(\fifo[13][6] ),
	.SE(n355),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[13][7] ),
	.D(n190),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[13][6]  (
	.SI(\fifo[13][5] ),
	.SE(n358),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[13][6] ),
	.D(n189),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[13][5]  (
	.SI(\fifo[13][4] ),
	.SE(n357),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[13][5] ),
	.D(n188),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[13][4]  (
	.SI(\fifo[13][3] ),
	.SE(n356),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[13][4] ),
	.D(n187),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[13][3]  (
	.SI(\fifo[13][2] ),
	.SE(n355),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[13][3] ),
	.D(n186),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[13][2]  (
	.SI(\fifo[13][1] ),
	.SE(n358),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[13][2] ),
	.D(n185),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[13][1]  (
	.SI(\fifo[13][0] ),
	.SE(n357),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[13][1] ),
	.D(n184),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[13][0]  (
	.SI(\fifo[12][7] ),
	.SE(n356),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[13][0] ),
	.D(n183),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[3][7]  (
	.SI(\fifo[3][6] ),
	.SE(n355),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[3][7] ),
	.D(n270),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[3][6]  (
	.SI(\fifo[3][5] ),
	.SE(n358),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[3][6] ),
	.D(n269),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[3][5]  (
	.SI(\fifo[3][4] ),
	.SE(n357),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[3][5] ),
	.D(n268),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[3][4]  (
	.SI(\fifo[3][3] ),
	.SE(n356),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[3][4] ),
	.D(n267),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[3][3]  (
	.SI(\fifo[3][2] ),
	.SE(n355),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[3][3] ),
	.D(n266),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[3][2]  (
	.SI(\fifo[3][1] ),
	.SE(n358),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[3][2] ),
	.D(n265),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[3][1]  (
	.SI(\fifo[3][0] ),
	.SE(n357),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[3][1] ),
	.D(n264),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[3][0]  (
	.SI(\fifo[2][7] ),
	.SE(n356),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[3][0] ),
	.D(n263),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[7][7]  (
	.SI(\fifo[7][6] ),
	.SE(n355),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[7][7] ),
	.D(n238),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[7][6]  (
	.SI(\fifo[7][5] ),
	.SE(n358),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[7][6] ),
	.D(n237),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[7][5]  (
	.SI(\fifo[7][4] ),
	.SE(n357),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[7][5] ),
	.D(n236),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[7][4]  (
	.SI(\fifo[7][3] ),
	.SE(n356),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[7][4] ),
	.D(n235),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[7][3]  (
	.SI(\fifo[7][2] ),
	.SE(n355),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[7][3] ),
	.D(n234),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[7][2]  (
	.SI(\fifo[7][1] ),
	.SE(n358),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[7][2] ),
	.D(n233),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[7][1]  (
	.SI(\fifo[7][0] ),
	.SE(n357),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[7][1] ),
	.D(n232),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[7][0]  (
	.SI(\fifo[6][7] ),
	.SE(n356),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[7][0] ),
	.D(n231),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[11][7]  (
	.SI(\fifo[11][6] ),
	.SE(n355),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[11][7] ),
	.D(n206),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[11][6]  (
	.SI(\fifo[11][5] ),
	.SE(n358),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[11][6] ),
	.D(n205),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[11][5]  (
	.SI(\fifo[11][4] ),
	.SE(n357),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[11][5] ),
	.D(n204),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[11][4]  (
	.SI(\fifo[11][3] ),
	.SE(n356),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[11][4] ),
	.D(n203),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[11][3]  (
	.SI(\fifo[11][2] ),
	.SE(n355),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[11][3] ),
	.D(n202),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[11][2]  (
	.SI(\fifo[11][1] ),
	.SE(n358),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[11][2] ),
	.D(n201),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[11][1]  (
	.SI(\fifo[11][0] ),
	.SE(n357),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[11][1] ),
	.D(n200),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[11][0]  (
	.SI(\fifo[10][7] ),
	.SE(n356),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[11][0] ),
	.D(n199),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[15][7]  (
	.SI(\fifo[15][6] ),
	.SE(n355),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[15][7] ),
	.D(n174),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[15][6]  (
	.SI(\fifo[15][5] ),
	.SE(n358),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[15][6] ),
	.D(n173),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[15][5]  (
	.SI(\fifo[15][4] ),
	.SE(n357),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[15][5] ),
	.D(n172),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[15][4]  (
	.SI(\fifo[15][3] ),
	.SE(n356),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[15][4] ),
	.D(n171),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[15][3]  (
	.SI(test_si3),
	.SE(n355),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[15][3] ),
	.D(n170),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[15][1]  (
	.SI(\fifo[15][0] ),
	.SE(n357),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[15][1] ),
	.D(n168),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[15][0]  (
	.SI(\fifo[14][7] ),
	.SE(n356),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[15][0] ),
	.D(n167),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[2][7]  (
	.SI(\fifo[2][6] ),
	.SE(n355),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[2][7] ),
	.D(n278),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[2][6]  (
	.SI(\fifo[2][5] ),
	.SE(n358),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[2][6] ),
	.D(n277),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[2][5]  (
	.SI(\fifo[2][4] ),
	.SE(n357),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[2][5] ),
	.D(n276),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[2][4]  (
	.SI(\fifo[2][3] ),
	.SE(n356),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[2][4] ),
	.D(n275),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[2][3]  (
	.SI(\fifo[2][2] ),
	.SE(n355),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[2][3] ),
	.D(n274),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[2][2]  (
	.SI(\fifo[2][1] ),
	.SE(n358),
	.RN(w_rst_n),
	.Q(\fifo[2][2] ),
	.D(n273),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[2][1]  (
	.SI(\fifo[2][0] ),
	.SE(n357),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[2][1] ),
	.D(n272),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[2][0]  (
	.SI(\fifo[1][7] ),
	.SE(n356),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[2][0] ),
	.D(n271),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[6][7]  (
	.SI(\fifo[6][6] ),
	.SE(n355),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[6][7] ),
	.D(n246),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[6][6]  (
	.SI(\fifo[6][5] ),
	.SE(n358),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[6][6] ),
	.D(n245),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[6][5]  (
	.SI(\fifo[6][4] ),
	.SE(n357),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[6][5] ),
	.D(n244),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[6][4]  (
	.SI(\fifo[6][3] ),
	.SE(n356),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[6][4] ),
	.D(n243),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[6][3]  (
	.SI(\fifo[6][2] ),
	.SE(n355),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[6][3] ),
	.D(n242),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[6][2]  (
	.SI(\fifo[6][1] ),
	.SE(n358),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[6][2] ),
	.D(n241),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[6][1]  (
	.SI(\fifo[6][0] ),
	.SE(n357),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[6][1] ),
	.D(n240),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[6][0]  (
	.SI(\fifo[5][7] ),
	.SE(n356),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[6][0] ),
	.D(n239),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[10][7]  (
	.SI(\fifo[10][6] ),
	.SE(n355),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[10][7] ),
	.D(n214),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[10][6]  (
	.SI(\fifo[10][5] ),
	.SE(n358),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[10][6] ),
	.D(n213),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[10][5]  (
	.SI(\fifo[10][4] ),
	.SE(n357),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[10][5] ),
	.D(n212),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[10][4]  (
	.SI(\fifo[10][3] ),
	.SE(n356),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[10][4] ),
	.D(n211),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[10][3]  (
	.SI(\fifo[10][2] ),
	.SE(n355),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[10][3] ),
	.D(n210),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[10][2]  (
	.SI(\fifo[10][1] ),
	.SE(n358),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[10][2] ),
	.D(n209),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[10][1]  (
	.SI(\fifo[10][0] ),
	.SE(n357),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[10][1] ),
	.D(n208),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[10][0]  (
	.SI(\fifo[9][7] ),
	.SE(n356),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[10][0] ),
	.D(n207),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[14][7]  (
	.SI(\fifo[14][6] ),
	.SE(n355),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[14][7] ),
	.D(n182),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[14][6]  (
	.SI(\fifo[14][5] ),
	.SE(n358),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[14][6] ),
	.D(n181),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[14][5]  (
	.SI(\fifo[14][4] ),
	.SE(n357),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[14][5] ),
	.D(n180),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[14][4]  (
	.SI(\fifo[14][3] ),
	.SE(n356),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[14][4] ),
	.D(n179),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[14][3]  (
	.SI(\fifo[14][2] ),
	.SE(n355),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[14][3] ),
	.D(n178),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[14][2]  (
	.SI(\fifo[14][1] ),
	.SE(n358),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[14][2] ),
	.D(n177),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[14][1]  (
	.SI(\fifo[14][0] ),
	.SE(n357),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[14][1] ),
	.D(n176),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[14][0]  (
	.SI(\fifo[13][7] ),
	.SE(n356),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[14][0] ),
	.D(n175),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[0][7]  (
	.SI(\fifo[0][6] ),
	.SE(n355),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[0][7] ),
	.D(n294),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[0][6]  (
	.SI(\fifo[0][5] ),
	.SE(n358),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[0][6] ),
	.D(n293),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[0][5]  (
	.SI(\fifo[0][4] ),
	.SE(n357),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[0][5] ),
	.D(n292),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[0][4]  (
	.SI(\fifo[0][3] ),
	.SE(n356),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[0][4] ),
	.D(n291),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[0][3]  (
	.SI(\fifo[0][2] ),
	.SE(n355),
	.RN(w_rst_n),
	.Q(\fifo[0][3] ),
	.D(n290),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[0][2]  (
	.SI(\fifo[0][1] ),
	.SE(n358),
	.RN(w_rst_n),
	.Q(\fifo[0][2] ),
	.D(n289),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[0][1]  (
	.SI(\fifo[0][0] ),
	.SE(n357),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[0][1] ),
	.D(n288),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[0][0]  (
	.SI(test_si1),
	.SE(n356),
	.RN(w_rst_n),
	.Q(\fifo[0][0] ),
	.D(n287),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[4][7]  (
	.SI(\fifo[4][6] ),
	.SE(n355),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[4][7] ),
	.D(n262),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[4][6]  (
	.SI(\fifo[4][5] ),
	.SE(n358),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[4][6] ),
	.D(n261),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[4][5]  (
	.SI(\fifo[4][4] ),
	.SE(n357),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[4][5] ),
	.D(n260),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[4][4]  (
	.SI(\fifo[4][3] ),
	.SE(n356),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[4][4] ),
	.D(n259),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[4][3]  (
	.SI(\fifo[4][2] ),
	.SE(n355),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[4][3] ),
	.D(n258),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[4][2]  (
	.SI(\fifo[4][1] ),
	.SE(n358),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[4][2] ),
	.D(n257),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[4][1]  (
	.SI(\fifo[4][0] ),
	.SE(n357),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[4][1] ),
	.D(n256),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[4][0]  (
	.SI(\fifo[3][7] ),
	.SE(n356),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[4][0] ),
	.D(n255),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[8][7]  (
	.SI(\fifo[8][6] ),
	.SE(n355),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[8][7] ),
	.D(n230),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[8][6]  (
	.SI(\fifo[8][5] ),
	.SE(n358),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[8][6] ),
	.D(n229),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[8][5]  (
	.SI(\fifo[8][4] ),
	.SE(n357),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[8][5] ),
	.D(n228),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[8][4]  (
	.SI(\fifo[8][3] ),
	.SE(n356),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[8][4] ),
	.D(n227),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[8][3]  (
	.SI(\fifo[8][2] ),
	.SE(n355),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[8][3] ),
	.D(n226),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[8][2]  (
	.SI(\fifo[8][1] ),
	.SE(n358),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[8][2] ),
	.D(n225),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[8][1]  (
	.SI(\fifo[8][0] ),
	.SE(n357),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[8][1] ),
	.D(n224),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[8][0]  (
	.SI(\fifo[7][7] ),
	.SE(n356),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[8][0] ),
	.D(n223),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[12][7]  (
	.SI(\fifo[12][6] ),
	.SE(n355),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[12][7] ),
	.D(n198),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[12][6]  (
	.SI(\fifo[12][5] ),
	.SE(n358),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[12][6] ),
	.D(n197),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[12][5]  (
	.SI(\fifo[12][4] ),
	.SE(n357),
	.RN(FE_OFN4_scan_rst_sync1_mux_out),
	.Q(\fifo[12][5] ),
	.D(n196),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[12][4]  (
	.SI(\fifo[12][3] ),
	.SE(n356),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[12][4] ),
	.D(n195),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[12][3]  (
	.SI(\fifo[12][2] ),
	.SE(n355),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[12][3] ),
	.D(n194),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[12][2]  (
	.SI(\fifo[12][1] ),
	.SE(n358),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[12][2] ),
	.D(n193),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[12][1]  (
	.SI(\fifo[12][0] ),
	.SE(n357),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[12][1] ),
	.D(n192),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \fifo_reg[12][0]  (
	.SI(\fifo[11][7] ),
	.SE(n356),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(\fifo[12][0] ),
	.D(n191),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U130 (
	.Y(n141),
	.B(n341),
	.A(n342), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U131 (
	.Y(n152),
	.B(w_address[2]),
	.A(w_address[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U132 (
	.Y(n146),
	.B(w_address[1]),
	.A(n342), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U133 (
	.Y(n149),
	.B(w_address[2]),
	.A(n341), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U149 (
	.Y(n143),
	.B(n141),
	.A(n144), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U150 (
	.Y(n158),
	.B(n141),
	.A(n159), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U151 (
	.Y(n322),
	.A(n319), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U152 (
	.Y(n321),
	.A(n319), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U153 (
	.Y(n318),
	.A(n316), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U156 (
	.Y(n145),
	.B(n142),
	.A(n146), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U157 (
	.Y(n147),
	.B(n144),
	.A(n146), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U158 (
	.Y(n148),
	.B(n142),
	.A(n149), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U159 (
	.Y(n150),
	.B(n144),
	.A(n149), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U160 (
	.Y(n151),
	.B(n142),
	.A(n152), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U161 (
	.Y(n154),
	.B(n144),
	.A(n152), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U162 (
	.Y(n160),
	.B(n146),
	.A(n157), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U163 (
	.Y(n161),
	.B(n146),
	.A(n159), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U164 (
	.Y(n162),
	.B(n149),
	.A(n157), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U165 (
	.Y(n163),
	.B(n149),
	.A(n159), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U166 (
	.Y(n164),
	.B(n152),
	.A(n157), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U167 (
	.Y(n166),
	.B(n152),
	.A(n159), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U168 (
	.Y(n156),
	.B(n141),
	.A(n157), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U169 (
	.Y(n140),
	.B(n142),
	.A(n141), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U170 (
	.Y(n144),
	.B(n340),
	.A(n153), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U171 (
	.Y(n155),
	.B(full_flag),
	.AN(w_inc), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U172 (
	.Y(n159),
	.B(n340),
	.A(n165), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U175 (
	.Y(n343),
	.A(w_data[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U176 (
	.Y(n344),
	.A(w_data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U177 (
	.Y(n345),
	.A(w_data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U178 (
	.Y(n346),
	.A(w_data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U179 (
	.Y(n347),
	.A(w_data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U180 (
	.Y(n348),
	.A(w_data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U181 (
	.Y(n349),
	.A(w_data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U182 (
	.Y(n350),
	.A(w_data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U183 (
	.Y(rd_data[6]),
	.S1(N11),
	.S0(N12),
	.D(n308),
	.C(n310),
	.B(n309),
	.A(n311), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U184 (
	.Y(n311),
	.S1(N10),
	.S0(n321),
	.D(\fifo[3][6] ),
	.C(\fifo[2][6] ),
	.B(\fifo[1][6] ),
	.A(\fifo[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U185 (
	.Y(n309),
	.S1(N10),
	.S0(n321),
	.D(\fifo[11][6] ),
	.C(\fifo[10][6] ),
	.B(\fifo[9][6] ),
	.A(\fifo[8][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U186 (
	.Y(n310),
	.S1(N10),
	.S0(n321),
	.D(\fifo[7][6] ),
	.C(\fifo[6][6] ),
	.B(\fifo[5][6] ),
	.A(\fifo[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U187 (
	.Y(rd_data[7]),
	.S1(N11),
	.S0(N12),
	.D(n312),
	.C(n314),
	.B(n313),
	.A(n315), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U188 (
	.Y(n315),
	.S1(N10),
	.S0(N9),
	.D(\fifo[3][7] ),
	.C(\fifo[2][7] ),
	.B(\fifo[1][7] ),
	.A(\fifo[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U189 (
	.Y(n313),
	.S1(N10),
	.S0(N9),
	.D(\fifo[11][7] ),
	.C(\fifo[10][7] ),
	.B(\fifo[9][7] ),
	.A(\fifo[8][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U190 (
	.Y(n314),
	.S1(N10),
	.S0(N9),
	.D(\fifo[7][7] ),
	.C(\fifo[6][7] ),
	.B(\fifo[5][7] ),
	.A(\fifo[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U191 (
	.Y(rd_data[2]),
	.S1(N11),
	.S0(N12),
	.D(n137),
	.C(n139),
	.B(n138),
	.A(n295), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U192 (
	.Y(n295),
	.S1(n318),
	.S0(n322),
	.D(\fifo[3][2] ),
	.C(\fifo[2][2] ),
	.B(\fifo[1][2] ),
	.A(\fifo[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U193 (
	.Y(n138),
	.S1(n318),
	.S0(n322),
	.D(\fifo[11][2] ),
	.C(\fifo[10][2] ),
	.B(\fifo[9][2] ),
	.A(\fifo[8][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U194 (
	.Y(n139),
	.S1(n318),
	.S0(n322),
	.D(\fifo[7][2] ),
	.C(\fifo[6][2] ),
	.B(\fifo[5][2] ),
	.A(\fifo[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U195 (
	.Y(n167),
	.B1(n343),
	.B0(n140),
	.A1N(n140),
	.A0N(\fifo[15][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U196 (
	.Y(n168),
	.B1(n344),
	.B0(n140),
	.A1N(n140),
	.A0N(\fifo[15][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U197 (
	.Y(n169),
	.B1(n345),
	.B0(n140),
	.A1N(n140),
	.A0N(n362), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U198 (
	.Y(n170),
	.B1(n346),
	.B0(n140),
	.A1N(n140),
	.A0N(\fifo[15][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U199 (
	.Y(n171),
	.B1(n347),
	.B0(n140),
	.A1N(n140),
	.A0N(\fifo[15][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U200 (
	.Y(n172),
	.B1(n348),
	.B0(n140),
	.A1N(n140),
	.A0N(\fifo[15][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U201 (
	.Y(n173),
	.B1(n349),
	.B0(n140),
	.A1N(n140),
	.A0N(\fifo[15][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U202 (
	.Y(n174),
	.B1(n350),
	.B0(n140),
	.A1N(n140),
	.A0N(\fifo[15][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U203 (
	.Y(n183),
	.B1(n145),
	.B0(n343),
	.A1N(n145),
	.A0N(\fifo[13][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U204 (
	.Y(n184),
	.B1(n145),
	.B0(n344),
	.A1N(n145),
	.A0N(\fifo[13][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U205 (
	.Y(n185),
	.B1(n145),
	.B0(n345),
	.A1N(n145),
	.A0N(\fifo[13][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U206 (
	.Y(n186),
	.B1(n145),
	.B0(n346),
	.A1N(n145),
	.A0N(\fifo[13][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U207 (
	.Y(n187),
	.B1(n145),
	.B0(n347),
	.A1N(n145),
	.A0N(\fifo[13][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U208 (
	.Y(n188),
	.B1(n145),
	.B0(n348),
	.A1N(n145),
	.A0N(\fifo[13][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U209 (
	.Y(n189),
	.B1(n145),
	.B0(n349),
	.A1N(n145),
	.A0N(\fifo[13][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U210 (
	.Y(n190),
	.B1(n145),
	.B0(n350),
	.A1N(n145),
	.A0N(\fifo[13][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U211 (
	.Y(n191),
	.B1(n147),
	.B0(n343),
	.A1N(n147),
	.A0N(\fifo[12][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U212 (
	.Y(n192),
	.B1(n147),
	.B0(n344),
	.A1N(n147),
	.A0N(\fifo[12][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U213 (
	.Y(n193),
	.B1(n147),
	.B0(n345),
	.A1N(n147),
	.A0N(\fifo[12][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U214 (
	.Y(n194),
	.B1(n147),
	.B0(n346),
	.A1N(n147),
	.A0N(\fifo[12][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U215 (
	.Y(n195),
	.B1(n147),
	.B0(n347),
	.A1N(n147),
	.A0N(\fifo[12][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U216 (
	.Y(n196),
	.B1(n147),
	.B0(n348),
	.A1N(n147),
	.A0N(\fifo[12][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U217 (
	.Y(n197),
	.B1(n147),
	.B0(n349),
	.A1N(n147),
	.A0N(\fifo[12][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U218 (
	.Y(n198),
	.B1(n147),
	.B0(n350),
	.A1N(n147),
	.A0N(\fifo[12][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U219 (
	.Y(n199),
	.B1(n148),
	.B0(n343),
	.A1N(n148),
	.A0N(\fifo[11][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U220 (
	.Y(n200),
	.B1(n148),
	.B0(n344),
	.A1N(n148),
	.A0N(\fifo[11][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U221 (
	.Y(n201),
	.B1(n148),
	.B0(n345),
	.A1N(n148),
	.A0N(\fifo[11][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U222 (
	.Y(n202),
	.B1(n148),
	.B0(n346),
	.A1N(n148),
	.A0N(\fifo[11][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U223 (
	.Y(n203),
	.B1(n148),
	.B0(n347),
	.A1N(n148),
	.A0N(\fifo[11][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U224 (
	.Y(n204),
	.B1(n148),
	.B0(n348),
	.A1N(n148),
	.A0N(\fifo[11][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U225 (
	.Y(n205),
	.B1(n148),
	.B0(n349),
	.A1N(n148),
	.A0N(\fifo[11][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U226 (
	.Y(n206),
	.B1(n148),
	.B0(n350),
	.A1N(n148),
	.A0N(\fifo[11][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U227 (
	.Y(n207),
	.B1(n150),
	.B0(n343),
	.A1N(n150),
	.A0N(\fifo[10][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U228 (
	.Y(n208),
	.B1(n150),
	.B0(n344),
	.A1N(n150),
	.A0N(\fifo[10][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U229 (
	.Y(n209),
	.B1(n150),
	.B0(n345),
	.A1N(n150),
	.A0N(\fifo[10][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U230 (
	.Y(n210),
	.B1(n150),
	.B0(n346),
	.A1N(n150),
	.A0N(\fifo[10][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U231 (
	.Y(n211),
	.B1(n150),
	.B0(n347),
	.A1N(n150),
	.A0N(\fifo[10][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U232 (
	.Y(n212),
	.B1(n150),
	.B0(n348),
	.A1N(n150),
	.A0N(\fifo[10][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U233 (
	.Y(n213),
	.B1(n150),
	.B0(n349),
	.A1N(n150),
	.A0N(\fifo[10][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U234 (
	.Y(n214),
	.B1(n150),
	.B0(n350),
	.A1N(n150),
	.A0N(\fifo[10][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U235 (
	.Y(n215),
	.B1(n151),
	.B0(n343),
	.A1N(n151),
	.A0N(\fifo[9][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U236 (
	.Y(n216),
	.B1(n151),
	.B0(n344),
	.A1N(n151),
	.A0N(\fifo[9][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U237 (
	.Y(n217),
	.B1(n151),
	.B0(n345),
	.A1N(n151),
	.A0N(\fifo[9][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U238 (
	.Y(n218),
	.B1(n151),
	.B0(n346),
	.A1N(n151),
	.A0N(\fifo[9][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U239 (
	.Y(n219),
	.B1(n151),
	.B0(n347),
	.A1N(n151),
	.A0N(\fifo[9][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U240 (
	.Y(n220),
	.B1(n151),
	.B0(n348),
	.A1N(n151),
	.A0N(\fifo[9][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U241 (
	.Y(n221),
	.B1(n151),
	.B0(n349),
	.A1N(n151),
	.A0N(\fifo[9][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U242 (
	.Y(n222),
	.B1(n151),
	.B0(n350),
	.A1N(n151),
	.A0N(\fifo[9][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U243 (
	.Y(n223),
	.B1(n154),
	.B0(n343),
	.A1N(n154),
	.A0N(\fifo[8][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U244 (
	.Y(n224),
	.B1(n154),
	.B0(n344),
	.A1N(n154),
	.A0N(\fifo[8][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U245 (
	.Y(n225),
	.B1(n154),
	.B0(n345),
	.A1N(n154),
	.A0N(\fifo[8][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U246 (
	.Y(n226),
	.B1(n154),
	.B0(n346),
	.A1N(n154),
	.A0N(\fifo[8][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U247 (
	.Y(n227),
	.B1(n154),
	.B0(n347),
	.A1N(n154),
	.A0N(\fifo[8][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U248 (
	.Y(n228),
	.B1(n154),
	.B0(n348),
	.A1N(n154),
	.A0N(\fifo[8][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U249 (
	.Y(n229),
	.B1(n154),
	.B0(n349),
	.A1N(n154),
	.A0N(\fifo[8][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U250 (
	.Y(n230),
	.B1(n154),
	.B0(n350),
	.A1N(n154),
	.A0N(\fifo[8][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U251 (
	.Y(n175),
	.B1(n143),
	.B0(n343),
	.A1N(n143),
	.A0N(\fifo[14][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U252 (
	.Y(n176),
	.B1(n143),
	.B0(n344),
	.A1N(n143),
	.A0N(\fifo[14][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U253 (
	.Y(n177),
	.B1(n143),
	.B0(n345),
	.A1N(n143),
	.A0N(\fifo[14][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U254 (
	.Y(n178),
	.B1(n143),
	.B0(n346),
	.A1N(n143),
	.A0N(\fifo[14][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U255 (
	.Y(n179),
	.B1(n143),
	.B0(n347),
	.A1N(n143),
	.A0N(\fifo[14][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U256 (
	.Y(n180),
	.B1(n143),
	.B0(n348),
	.A1N(n143),
	.A0N(\fifo[14][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U257 (
	.Y(n181),
	.B1(n143),
	.B0(n349),
	.A1N(n143),
	.A0N(\fifo[14][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U258 (
	.Y(n182),
	.B1(n143),
	.B0(n350),
	.A1N(n143),
	.A0N(\fifo[14][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U259 (
	.Y(n231),
	.B1(n156),
	.B0(n343),
	.A1N(n156),
	.A0N(\fifo[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U260 (
	.Y(n232),
	.B1(n156),
	.B0(n344),
	.A1N(n156),
	.A0N(\fifo[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U261 (
	.Y(n233),
	.B1(n156),
	.B0(n345),
	.A1N(n156),
	.A0N(\fifo[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U262 (
	.Y(n234),
	.B1(n156),
	.B0(n346),
	.A1N(n156),
	.A0N(\fifo[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U263 (
	.Y(n235),
	.B1(n156),
	.B0(n347),
	.A1N(n156),
	.A0N(\fifo[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U264 (
	.Y(n236),
	.B1(n156),
	.B0(n348),
	.A1N(n156),
	.A0N(\fifo[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U265 (
	.Y(n237),
	.B1(n156),
	.B0(n349),
	.A1N(n156),
	.A0N(\fifo[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U266 (
	.Y(n238),
	.B1(n156),
	.B0(n350),
	.A1N(n156),
	.A0N(\fifo[7][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U267 (
	.Y(n239),
	.B1(n158),
	.B0(n343),
	.A1N(n158),
	.A0N(\fifo[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U268 (
	.Y(n240),
	.B1(n158),
	.B0(n344),
	.A1N(n158),
	.A0N(\fifo[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U269 (
	.Y(n241),
	.B1(n158),
	.B0(n345),
	.A1N(n158),
	.A0N(\fifo[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U270 (
	.Y(n242),
	.B1(n158),
	.B0(n346),
	.A1N(n158),
	.A0N(\fifo[6][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U271 (
	.Y(n243),
	.B1(n158),
	.B0(n347),
	.A1N(n158),
	.A0N(\fifo[6][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U272 (
	.Y(n244),
	.B1(n158),
	.B0(n348),
	.A1N(n158),
	.A0N(\fifo[6][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U273 (
	.Y(n245),
	.B1(n158),
	.B0(n349),
	.A1N(n158),
	.A0N(\fifo[6][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U274 (
	.Y(n246),
	.B1(n158),
	.B0(n350),
	.A1N(n158),
	.A0N(\fifo[6][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U275 (
	.Y(n247),
	.B1(n160),
	.B0(n343),
	.A1N(n160),
	.A0N(n360), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U276 (
	.Y(n248),
	.B1(n160),
	.B0(n344),
	.A1N(n160),
	.A0N(\fifo[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U277 (
	.Y(n249),
	.B1(n160),
	.B0(n345),
	.A1N(n160),
	.A0N(\fifo[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U278 (
	.Y(n250),
	.B1(n160),
	.B0(n346),
	.A1N(n160),
	.A0N(\fifo[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U279 (
	.Y(n251),
	.B1(n160),
	.B0(n347),
	.A1N(n160),
	.A0N(\fifo[5][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U280 (
	.Y(n252),
	.B1(n160),
	.B0(n348),
	.A1N(n160),
	.A0N(\fifo[5][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U281 (
	.Y(n253),
	.B1(n160),
	.B0(n349),
	.A1N(n160),
	.A0N(\fifo[5][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U282 (
	.Y(n254),
	.B1(n160),
	.B0(n350),
	.A1N(n160),
	.A0N(\fifo[5][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U283 (
	.Y(n255),
	.B1(n161),
	.B0(n343),
	.A1N(n161),
	.A0N(\fifo[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U284 (
	.Y(n256),
	.B1(n161),
	.B0(n344),
	.A1N(n161),
	.A0N(\fifo[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U285 (
	.Y(n257),
	.B1(n161),
	.B0(n345),
	.A1N(n161),
	.A0N(\fifo[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U286 (
	.Y(n258),
	.B1(n161),
	.B0(n346),
	.A1N(n161),
	.A0N(\fifo[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U287 (
	.Y(n259),
	.B1(n161),
	.B0(n347),
	.A1N(n161),
	.A0N(\fifo[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U288 (
	.Y(n260),
	.B1(n161),
	.B0(n348),
	.A1N(n161),
	.A0N(\fifo[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U289 (
	.Y(n261),
	.B1(n161),
	.B0(n349),
	.A1N(n161),
	.A0N(\fifo[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U290 (
	.Y(n262),
	.B1(n161),
	.B0(n350),
	.A1N(n161),
	.A0N(\fifo[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U291 (
	.Y(n263),
	.B1(n162),
	.B0(n343),
	.A1N(n162),
	.A0N(\fifo[3][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U292 (
	.Y(n264),
	.B1(n162),
	.B0(n344),
	.A1N(n162),
	.A0N(\fifo[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U293 (
	.Y(n265),
	.B1(n162),
	.B0(n345),
	.A1N(n162),
	.A0N(\fifo[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U294 (
	.Y(n266),
	.B1(n162),
	.B0(n346),
	.A1N(n162),
	.A0N(\fifo[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U295 (
	.Y(n267),
	.B1(n162),
	.B0(n347),
	.A1N(n162),
	.A0N(\fifo[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U296 (
	.Y(n268),
	.B1(n162),
	.B0(n348),
	.A1N(n162),
	.A0N(\fifo[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U297 (
	.Y(n269),
	.B1(n162),
	.B0(n349),
	.A1N(n162),
	.A0N(\fifo[3][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U298 (
	.Y(n270),
	.B1(n162),
	.B0(n350),
	.A1N(n162),
	.A0N(\fifo[3][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U299 (
	.Y(n271),
	.B1(n163),
	.B0(n343),
	.A1N(n163),
	.A0N(\fifo[2][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U300 (
	.Y(n272),
	.B1(n163),
	.B0(n344),
	.A1N(n163),
	.A0N(\fifo[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U301 (
	.Y(n273),
	.B1(n163),
	.B0(n345),
	.A1N(n163),
	.A0N(\fifo[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U302 (
	.Y(n274),
	.B1(n163),
	.B0(n346),
	.A1N(n163),
	.A0N(\fifo[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U303 (
	.Y(n275),
	.B1(n163),
	.B0(n347),
	.A1N(n163),
	.A0N(\fifo[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U304 (
	.Y(n276),
	.B1(n163),
	.B0(n348),
	.A1N(n163),
	.A0N(\fifo[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U305 (
	.Y(n277),
	.B1(n163),
	.B0(n349),
	.A1N(n163),
	.A0N(\fifo[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U306 (
	.Y(n278),
	.B1(n163),
	.B0(n350),
	.A1N(n163),
	.A0N(\fifo[2][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U307 (
	.Y(n279),
	.B1(n164),
	.B0(n343),
	.A1N(n164),
	.A0N(\fifo[1][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U308 (
	.Y(n280),
	.B1(n164),
	.B0(n344),
	.A1N(n164),
	.A0N(\fifo[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U309 (
	.Y(n281),
	.B1(n164),
	.B0(n345),
	.A1N(n164),
	.A0N(\fifo[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U310 (
	.Y(n282),
	.B1(n164),
	.B0(n346),
	.A1N(n164),
	.A0N(\fifo[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U311 (
	.Y(n283),
	.B1(n164),
	.B0(n347),
	.A1N(n164),
	.A0N(\fifo[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U312 (
	.Y(n284),
	.B1(n164),
	.B0(n348),
	.A1N(n164),
	.A0N(\fifo[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U313 (
	.Y(n285),
	.B1(n164),
	.B0(n349),
	.A1N(n164),
	.A0N(\fifo[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U314 (
	.Y(n286),
	.B1(n164),
	.B0(n350),
	.A1N(n164),
	.A0N(\fifo[1][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U315 (
	.Y(n287),
	.B1(n166),
	.B0(n343),
	.A1N(n166),
	.A0N(\fifo[0][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U316 (
	.Y(n288),
	.B1(n166),
	.B0(n344),
	.A1N(n166),
	.A0N(\fifo[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U317 (
	.Y(n289),
	.B1(n166),
	.B0(n345),
	.A1N(n166),
	.A0N(\fifo[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U318 (
	.Y(n290),
	.B1(n166),
	.B0(n346),
	.A1N(n166),
	.A0N(\fifo[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U319 (
	.Y(n291),
	.B1(n166),
	.B0(n347),
	.A1N(n166),
	.A0N(\fifo[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U320 (
	.Y(n292),
	.B1(n166),
	.B0(n348),
	.A1N(n166),
	.A0N(\fifo[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U321 (
	.Y(n293),
	.B1(n166),
	.B0(n349),
	.A1N(n166),
	.A0N(\fifo[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U322 (
	.Y(n294),
	.B1(n166),
	.B0(n350),
	.A1N(n166),
	.A0N(\fifo[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U323 (
	.Y(rd_data[3]),
	.S1(N11),
	.S0(N12),
	.D(n296),
	.C(n298),
	.B(n297),
	.A(n299), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U324 (
	.Y(n299),
	.S1(n318),
	.S0(n322),
	.D(\fifo[3][3] ),
	.C(\fifo[2][3] ),
	.B(\fifo[1][3] ),
	.A(\fifo[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U325 (
	.Y(n297),
	.S1(n318),
	.S0(n322),
	.D(\fifo[11][3] ),
	.C(\fifo[10][3] ),
	.B(\fifo[9][3] ),
	.A(\fifo[8][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U326 (
	.Y(n298),
	.S1(n318),
	.S0(n322),
	.D(\fifo[7][3] ),
	.C(\fifo[6][3] ),
	.B(\fifo[5][3] ),
	.A(\fifo[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U327 (
	.Y(n142),
	.B(w_address[0]),
	.A(n153), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U328 (
	.Y(n157),
	.B(w_address[0]),
	.A(n165), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U329 (
	.Y(n165),
	.B(w_address[3]),
	.AN(n155), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U330 (
	.Y(rd_data[4]),
	.S1(N11),
	.S0(N12),
	.D(n300),
	.C(n302),
	.B(n301),
	.A(n303), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U331 (
	.Y(n303),
	.S1(n318),
	.S0(n322),
	.D(\fifo[3][4] ),
	.C(\fifo[2][4] ),
	.B(\fifo[1][4] ),
	.A(\fifo[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U332 (
	.Y(n301),
	.S1(n318),
	.S0(n322),
	.D(\fifo[11][4] ),
	.C(\fifo[10][4] ),
	.B(\fifo[9][4] ),
	.A(\fifo[8][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U333 (
	.Y(n302),
	.S1(n318),
	.S0(n322),
	.D(\fifo[7][4] ),
	.C(\fifo[6][4] ),
	.B(\fifo[5][4] ),
	.A(\fifo[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U334 (
	.Y(rd_data[0]),
	.S1(N11),
	.S0(N12),
	.D(n129),
	.C(n131),
	.B(n130),
	.A(n132), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U335 (
	.Y(n132),
	.S1(N10),
	.S0(n321),
	.D(\fifo[3][0] ),
	.C(\fifo[2][0] ),
	.B(\fifo[1][0] ),
	.A(\fifo[0][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U336 (
	.Y(n130),
	.S1(N10),
	.S0(n321),
	.D(\fifo[11][0] ),
	.C(\fifo[10][0] ),
	.B(\fifo[9][0] ),
	.A(\fifo[8][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U337 (
	.Y(n131),
	.S1(N10),
	.S0(n321),
	.D(\fifo[7][0] ),
	.C(\fifo[6][0] ),
	.B(n360),
	.A(\fifo[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U338 (
	.Y(rd_data[5]),
	.S1(N11),
	.S0(N12),
	.D(n304),
	.C(n306),
	.B(n305),
	.A(n307), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U339 (
	.Y(n307),
	.S1(N10),
	.S0(n321),
	.D(\fifo[3][5] ),
	.C(\fifo[2][5] ),
	.B(\fifo[1][5] ),
	.A(\fifo[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U340 (
	.Y(n305),
	.S1(N10),
	.S0(n321),
	.D(\fifo[11][5] ),
	.C(\fifo[10][5] ),
	.B(\fifo[9][5] ),
	.A(\fifo[8][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U341 (
	.Y(n306),
	.S1(N10),
	.S0(n321),
	.D(\fifo[7][5] ),
	.C(\fifo[6][5] ),
	.B(\fifo[5][5] ),
	.A(\fifo[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U342 (
	.Y(rd_data[1]),
	.S1(N11),
	.S0(N12),
	.D(n133),
	.C(n135),
	.B(n134),
	.A(n136), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U343 (
	.Y(n134),
	.S1(N10),
	.S0(n321),
	.D(\fifo[11][1] ),
	.C(\fifo[10][1] ),
	.B(\fifo[9][1] ),
	.A(\fifo[8][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U344 (
	.Y(n133),
	.S1(n318),
	.S0(n321),
	.D(\fifo[15][1] ),
	.C(\fifo[14][1] ),
	.B(\fifo[13][1] ),
	.A(\fifo[12][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U345 (
	.Y(n136),
	.S1(N10),
	.S0(n322),
	.D(\fifo[3][1] ),
	.C(\fifo[2][1] ),
	.B(\fifo[1][1] ),
	.A(\fifo[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U346 (
	.Y(n135),
	.S1(N10),
	.S0(n322),
	.D(\fifo[7][1] ),
	.C(\fifo[6][1] ),
	.B(\fifo[5][1] ),
	.A(\fifo[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U347 (
	.Y(n129),
	.S1(N10),
	.S0(n321),
	.D(\fifo[15][0] ),
	.C(\fifo[14][0] ),
	.B(\fifo[13][0] ),
	.A(\fifo[12][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U348 (
	.Y(n308),
	.S1(N10),
	.S0(n321),
	.D(\fifo[15][6] ),
	.C(\fifo[14][6] ),
	.B(\fifo[13][6] ),
	.A(\fifo[12][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U349 (
	.Y(n312),
	.S1(N10),
	.S0(N9),
	.D(\fifo[15][7] ),
	.C(\fifo[14][7] ),
	.B(\fifo[13][7] ),
	.A(\fifo[12][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U350 (
	.Y(n137),
	.S1(n318),
	.S0(n322),
	.D(n362),
	.C(\fifo[14][2] ),
	.B(\fifo[13][2] ),
	.A(\fifo[12][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U351 (
	.Y(n296),
	.S1(n318),
	.S0(n322),
	.D(\fifo[15][3] ),
	.C(\fifo[14][3] ),
	.B(\fifo[13][3] ),
	.A(\fifo[12][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U352 (
	.Y(n300),
	.S1(n318),
	.S0(n322),
	.D(\fifo[15][4] ),
	.C(\fifo[14][4] ),
	.B(\fifo[13][4] ),
	.A(\fifo[12][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U353 (
	.Y(n304),
	.S1(n318),
	.S0(n321),
	.D(\fifo[15][5] ),
	.C(\fifo[14][5] ),
	.B(\fifo[13][5] ),
	.A(\fifo[12][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U354 (
	.Y(n153),
	.B(n155),
	.A(w_address[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U355 (
	.Y(n316),
	.A(N10), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U356 (
	.Y(n319),
	.A(N9), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U357 (
	.Y(n341),
	.A(w_address[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U358 (
	.Y(n342),
	.A(w_address[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U359 (
	.Y(n340),
	.A(w_address[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U360 (
	.Y(n355),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U361 (
	.Y(n356),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U362 (
	.Y(n357),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U363 (
	.Y(n358),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U364 (
	.Y(n359),
	.A(\fifo[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U365 (
	.Y(n360),
	.A(n359), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U366 (
	.Y(n361),
	.A(\fifo[15][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U367 (
	.Y(n362),
	.A(n361), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX4M \fifo_reg[5][0]  (
	.SI(\fifo[4][7] ),
	.SE(n356),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(FE_OFN9_SO_4_),
	.D(n247),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX4M \fifo_reg[15][2]  (
	.SI(\fifo[15][1] ),
	.SE(n358),
	.RN(FE_OFN3_scan_rst_sync1_mux_out),
	.Q(FE_OFN8_SO_3_),
	.D(n169),
	.CK(w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module empty_gen_test_1 (
	sync_grey_coded_wr_ptr, 
	rd_clk, 
	rd_rst_n, 
	rd_inc, 
	rd_ptr_grey_coded, 
	rd_address, 
	empty_flag, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input [4:0] sync_grey_coded_wr_ptr;
   input rd_clk;
   input rd_rst_n;
   input rd_inc;
   output [4:0] rd_ptr_grey_coded;
   output [3:0] rd_address;
   output empty_flag;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N7;
   wire N8;
   wire N9;
   wire N10;
   wire N11;
   wire n1;
   wire n3;
   wire n4;
   wire n5;
   wire n7;
   wire n9;
   wire n11;
   wire n13;
   wire n15;
   wire n17;
   wire n19;
   wire n21;
   wire n23;
   wire \add_23/carry[4] ;
   wire \add_23/carry[3] ;
   wire \add_23/carry[2] ;
   wire n2;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire [4:0] rd_ptr;

   assign test_so = rd_ptr[4] ;

   // Module instantiations
   SDFFRQX2M \rd_ptr_reg[4]  (
	.SI(rd_ptr[3]),
	.SE(test_se),
	.RN(rd_rst_n),
	.Q(rd_ptr[4]),
	.D(n21),
	.CK(rd_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \rd_ptr_reg[0]  (
	.SI(rd_address[3]),
	.SE(test_se),
	.RN(rd_rst_n),
	.Q(rd_ptr[0]),
	.D(n23),
	.CK(rd_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \rd_address_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(rd_rst_n),
	.Q(rd_address[0]),
	.D(n19),
	.CK(rd_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX4M \rd_address_reg[1]  (
	.SI(rd_address[0]),
	.SE(test_se),
	.RN(rd_rst_n),
	.Q(rd_address[1]),
	.D(n17),
	.CK(rd_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \rd_address_reg[2]  (
	.SI(rd_address[1]),
	.SE(test_se),
	.RN(rd_rst_n),
	.Q(rd_address[2]),
	.D(n15),
	.CK(rd_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \rd_ptr_reg[1]  (
	.SI(N7),
	.SE(test_se),
	.RN(rd_rst_n),
	.Q(rd_ptr[1]),
	.D(n11),
	.CK(rd_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \rd_ptr_reg[2]  (
	.SI(rd_ptr[1]),
	.SE(test_se),
	.RN(rd_rst_n),
	.Q(rd_ptr[2]),
	.D(n9),
	.CK(rd_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \rd_ptr_reg[3]  (
	.SI(rd_ptr[2]),
	.SE(test_se),
	.RN(rd_rst_n),
	.Q(rd_ptr[3]),
	.D(n7),
	.CK(rd_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \rd_address_reg[3]  (
	.SI(rd_address[2]),
	.SE(test_se),
	.RN(rd_rst_n),
	.Q(rd_address[3]),
	.D(n13),
	.CK(rd_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(n31),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U4 (
	.Y(n1),
	.B(rd_inc),
	.AN(empty_flag), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U5 (
	.Y(n15),
	.B(n4),
	.A(rd_address[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U6 (
	.Y(n4),
	.B(n5),
	.A(rd_address[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U7 (
	.Y(n5),
	.B(n31),
	.A(rd_address[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U8 (
	.Y(n7),
	.B1(n31),
	.B0(N10),
	.A1(n1),
	.A0(rd_ptr[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U9 (
	.Y(n9),
	.B1(n31),
	.B0(N9),
	.A1(n1),
	.A0(rd_ptr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U10 (
	.Y(n11),
	.B1(n31),
	.B0(N8),
	.A1(n1),
	.A0(rd_ptr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U11 (
	.Y(n21),
	.B1(n31),
	.B0(N11),
	.A1(n1),
	.A0(rd_ptr[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U12 (
	.Y(n23),
	.B1(n31),
	.B0(N7),
	.A1(n1),
	.A0(rd_ptr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U13 (
	.Y(n13),
	.B(n3),
	.A(rd_address[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U14 (
	.Y(n3),
	.B(n4),
	.AN(rd_address[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U15 (
	.Y(n17),
	.B(n5),
	.A(rd_address[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U16 (
	.Y(n19),
	.B(n31),
	.A(rd_address[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U26 (
	.S(N8),
	.CO(\add_23/carry[2] ),
	.B(rd_ptr[0]),
	.A(rd_ptr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U27 (
	.S(N9),
	.CO(\add_23/carry[3] ),
	.B(\add_23/carry[2] ),
	.A(rd_ptr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U28 (
	.S(N10),
	.CO(\add_23/carry[4] ),
	.B(\add_23/carry[3] ),
	.A(rd_ptr[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U29 (
	.Y(N7),
	.A(rd_ptr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U30 (
	.Y(N11),
	.B(rd_ptr[4]),
	.A(\add_23/carry[4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U31 (
	.Y(n30),
	.B(rd_ptr_grey_coded[2]),
	.A(sync_grey_coded_wr_ptr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U32 (
	.Y(n2),
	.B(rd_ptr_grey_coded[0]),
	.AN(sync_grey_coded_wr_ptr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U33 (
	.Y(n26),
	.B1(n2),
	.B0(sync_grey_coded_wr_ptr[1]),
	.A1N(rd_ptr_grey_coded[1]),
	.A0(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U34 (
	.Y(n24),
	.B(sync_grey_coded_wr_ptr[0]),
	.AN(rd_ptr_grey_coded[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U35 (
	.Y(n25),
	.B1(n24),
	.B0(rd_ptr_grey_coded[1]),
	.A1N(sync_grey_coded_wr_ptr[1]),
	.A0(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U36 (
	.Y(n29),
	.B(n25),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U37 (
	.Y(n28),
	.B(rd_ptr_grey_coded[3]),
	.A(sync_grey_coded_wr_ptr[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U38 (
	.Y(n27),
	.B(rd_ptr_grey_coded[4]),
	.A(sync_grey_coded_wr_ptr[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U39 (
	.Y(empty_flag),
	.D(n27),
	.C(n28),
	.B(n29),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   grey_code_gen_1 rd_ptr_gc (
	.binary_data({ rd_ptr[4],
		rd_ptr[3],
		rd_ptr[2],
		rd_ptr[1],
		rd_ptr[0] }),
	.grey_coded_data({ rd_ptr_grey_coded[4],
		rd_ptr_grey_coded[3],
		rd_ptr_grey_coded[2],
		rd_ptr_grey_coded[1],
		rd_ptr_grey_coded[0] }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module grey_code_gen_1 (
	binary_data, 
	grey_coded_data, 
	VDD, 
	VSS);
   input [4:0] binary_data;
   output [4:0] grey_coded_data;
   inout VDD;
   inout VSS;

   // Module instantiations
   CLKXOR2X2M U1 (
	.Y(grey_coded_data[1]),
	.B(binary_data[1]),
	.A(binary_data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U2 (
	.Y(grey_coded_data[0]),
	.B(binary_data[0]),
	.A(binary_data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U3 (
	.Y(grey_coded_data[2]),
	.B(binary_data[2]),
	.A(binary_data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U4 (
	.Y(grey_coded_data[3]),
	.B(binary_data[3]),
	.A(binary_data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U5 (
	.Y(grey_coded_data[4]),
	.A(binary_data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module synchronizer_test_0 (
	d1, 
	clk, 
	rst_n, 
	q2, 
	test_si, 
	test_se, 
	scan_clk_ref_clk_mux_out__L4_N1, 
	VDD, 
	VSS);
   input [4:0] d1;
   input clk;
   input rst_n;
   output [4:0] q2;
   input test_si;
   input test_se;
   input scan_clk_ref_clk_mux_out__L4_N1;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [4:0] q1;

   // Module instantiations
   SDFFRQX2M \q2_reg[4]  (
	.SI(q2[3]),
	.SE(test_se),
	.RN(rst_n),
	.Q(q2[4]),
	.D(q1[4]),
	.CK(scan_clk_ref_clk_mux_out__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \q2_reg[3]  (
	.SI(q2[2]),
	.SE(test_se),
	.RN(rst_n),
	.Q(q2[3]),
	.D(q1[3]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \q2_reg[2]  (
	.SI(q2[1]),
	.SE(test_se),
	.RN(rst_n),
	.Q(q2[2]),
	.D(q1[2]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \q2_reg[1]  (
	.SI(q2[0]),
	.SE(test_se),
	.RN(rst_n),
	.Q(q2[1]),
	.D(q1[1]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \q2_reg[0]  (
	.SI(q1[4]),
	.SE(test_se),
	.RN(rst_n),
	.Q(q2[0]),
	.D(q1[0]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \q1_reg[4]  (
	.SI(q1[3]),
	.SE(test_se),
	.RN(rst_n),
	.Q(q1[4]),
	.D(d1[4]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \q1_reg[3]  (
	.SI(q1[2]),
	.SE(test_se),
	.RN(rst_n),
	.Q(q1[3]),
	.D(d1[3]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \q1_reg[2]  (
	.SI(q1[1]),
	.SE(test_se),
	.RN(rst_n),
	.Q(q1[2]),
	.D(d1[2]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \q1_reg[1]  (
	.SI(q1[0]),
	.SE(test_se),
	.RN(rst_n),
	.Q(q1[1]),
	.D(d1[1]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \q1_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(rst_n),
	.Q(q1[0]),
	.D(d1[0]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module synchronizer_test_1 (
	d1, 
	clk, 
	rst_n, 
	q2, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input [4:0] d1;
   input clk;
   input rst_n;
   output [4:0] q2;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [4:0] q1;

   // Module instantiations
   SDFFRQX2M \q2_reg[0]  (
	.SI(q1[4]),
	.SE(test_se),
	.RN(rst_n),
	.Q(q2[0]),
	.D(q1[0]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \q2_reg[1]  (
	.SI(q2[0]),
	.SE(test_se),
	.RN(rst_n),
	.Q(q2[1]),
	.D(q1[1]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \q2_reg[4]  (
	.SI(q2[3]),
	.SE(test_se),
	.RN(rst_n),
	.Q(q2[4]),
	.D(q1[4]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \q2_reg[3]  (
	.SI(q2[2]),
	.SE(test_se),
	.RN(rst_n),
	.Q(q2[3]),
	.D(q1[3]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \q2_reg[2]  (
	.SI(q2[1]),
	.SE(test_se),
	.RN(rst_n),
	.Q(q2[2]),
	.D(q1[2]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \q1_reg[4]  (
	.SI(q1[3]),
	.SE(test_se),
	.RN(rst_n),
	.Q(q1[4]),
	.D(d1[4]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \q1_reg[3]  (
	.SI(q1[2]),
	.SE(test_se),
	.RN(rst_n),
	.Q(q1[3]),
	.D(d1[3]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \q1_reg[2]  (
	.SI(q1[1]),
	.SE(test_se),
	.RN(rst_n),
	.Q(q1[2]),
	.D(d1[2]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \q1_reg[1]  (
	.SI(q1[0]),
	.SE(test_se),
	.RN(rst_n),
	.Q(q1[1]),
	.D(d1[1]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \q1_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(rst_n),
	.Q(q1[0]),
	.D(d1[0]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module UART_tx_TOP_MODULE_test_1 (
	p_data, 
	clk, 
	rst_n, 
	data_valid, 
	parity_type, 
	parity_enable, 
	tx_out, 
	busy, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input [7:0] p_data;
   input clk;
   input rst_n;
   input data_valid;
   input parity_type;
   input parity_enable;
   output tx_out;
   output busy;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire serilaizer_done;
   wire serilaizer_enable;
   wire serialized_data;
   wire parity_bit;
   wire n3;
   wire n4;
   wire [1:0] mux_sel;

   assign test_so = parity_bit ;

   // Module instantiations
   fsm_controller_test_1 uut0 (
	.data_valid(data_valid),
	.serilaizer_done(serilaizer_done),
	.parity_enable(parity_enable),
	.clk(clk),
	.rst_n(rst_n),
	.serilaizer_enable(serilaizer_enable),
	.busy(busy),
	.mux_sel({ mux_sel[1],
		mux_sel[0] }),
	.test_si(test_si),
	.test_so(n4),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   serilaizer_test_1 uut1 (
	.p_data({ p_data[7],
		p_data[6],
		p_data[5],
		p_data[4],
		p_data[3],
		p_data[2],
		p_data[1],
		p_data[0] }),
	.data_valid(data_valid),
	.serilaizer_enable(serilaizer_enable),
	.busy(busy),
	.clk(clk),
	.rst_n(rst_n),
	.serialized_data(serialized_data),
	.serilaizer_done(serilaizer_done),
	.test_si(n4),
	.test_so(n3),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   parity_calc_test_1 uut2 (
	.p_data({ p_data[7],
		p_data[6],
		p_data[5],
		p_data[4],
		p_data[3],
		p_data[2],
		p_data[1],
		p_data[0] }),
	.data_valid(data_valid),
	.busy(busy),
	.parity_type(parity_type),
	.clk(clk),
	.rst_n(rst_n),
	.parity_bit(parity_bit),
	.test_si(n3),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   mux uu3 (
	.mux_sel({ mux_sel[1],
		mux_sel[0] }),
	.parity_bit(parity_bit),
	.serialized_data(serialized_data),
	.tx_out(tx_out), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module fsm_controller_test_1 (
	data_valid, 
	serilaizer_done, 
	parity_enable, 
	clk, 
	rst_n, 
	serilaizer_enable, 
	busy, 
	mux_sel, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input data_valid;
   input serilaizer_done;
   input parity_enable;
   input clk;
   input rst_n;
   output serilaizer_enable;
   output busy;
   output [1:0] mux_sel;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n4;
   wire n5;
   wire n6;
   wire [2:0] current_state;

   assign test_so = current_state[2] ;

   // Module instantiations
   SDFFRQX2M \current_state_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(rst_n),
	.Q(current_state[0]),
	.D(n17),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[2]  (
	.SI(n5),
	.SE(test_se),
	.RN(rst_n),
	.Q(current_state[2]),
	.D(n16),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[1]  (
	.SI(current_state[0]),
	.SE(test_se),
	.RN(rst_n),
	.Q(current_state[1]),
	.D(n15),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX2M U6 (
	.Y(busy),
	.C(n12),
	.B(n8),
	.AN(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U7 (
	.Y(serilaizer_enable),
	.B(n8),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U8 (
	.Y(n16),
	.B0(n12),
	.A1(n8),
	.A0(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U9 (
	.Y(n11),
	.B0(n7),
	.A1(n6),
	.A0(serilaizer_done), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U10 (
	.Y(n7),
	.B(n4),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U11 (
	.Y(n12),
	.B(current_state[0]),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U12 (
	.Y(n8),
	.B(n12),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U13 (
	.Y(n4),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U14 (
	.Y(n15),
	.B1(n5),
	.B0(n9),
	.A2(current_state[1]),
	.A1(current_state[2]),
	.A0(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U15 (
	.Y(n9),
	.B(n10),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U16 (
	.Y(n10),
	.B0(current_state[0]),
	.A1(n6),
	.A0(serilaizer_done), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U17 (
	.Y(n17),
	.B0(n7),
	.A2(n14),
	.A1(n12),
	.A0(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U18 (
	.Y(n14),
	.B(n5),
	.A(data_valid), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U19 (
	.Y(n13),
	.C(parity_enable),
	.B(current_state[1]),
	.A(serilaizer_done), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n5),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U21 (
	.Y(n6),
	.A(parity_enable), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U22 (
	.Y(mux_sel[0]),
	.B1(current_state[0]),
	.B0(current_state[1]),
	.A1N(mux_sel[1]),
	.A0N(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U23 (
	.Y(mux_sel[1]),
	.B(current_state[2]),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module serilaizer_test_1 (
	p_data, 
	data_valid, 
	serilaizer_enable, 
	busy, 
	clk, 
	rst_n, 
	serialized_data, 
	serilaizer_done, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input [7:0] p_data;
   input data_valid;
   input serilaizer_enable;
   input busy;
   input clk;
   input rst_n;
   output serialized_data;
   output serilaizer_done;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \counter[0] ;
   wire N24;
   wire N25;
   wire N26;
   wire n12;
   wire n13;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n14;
   wire n35;
   wire n36;
   wire [7:1] parallel_data_reg;

   assign test_so = parallel_data_reg[7] ;

   // Module instantiations
   SDFFRQX2M \parallel_data_reg_reg[6]  (
	.SI(parallel_data_reg[5]),
	.SE(test_se),
	.RN(rst_n),
	.Q(parallel_data_reg[6]),
	.D(n28),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \parallel_data_reg_reg[5]  (
	.SI(parallel_data_reg[4]),
	.SE(test_se),
	.RN(rst_n),
	.Q(parallel_data_reg[5]),
	.D(n29),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \parallel_data_reg_reg[4]  (
	.SI(parallel_data_reg[3]),
	.SE(test_se),
	.RN(rst_n),
	.Q(parallel_data_reg[4]),
	.D(n30),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \parallel_data_reg_reg[3]  (
	.SI(parallel_data_reg[2]),
	.SE(test_se),
	.RN(rst_n),
	.Q(parallel_data_reg[3]),
	.D(n31),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \parallel_data_reg_reg[2]  (
	.SI(parallel_data_reg[1]),
	.SE(test_se),
	.RN(rst_n),
	.Q(parallel_data_reg[2]),
	.D(n32),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \parallel_data_reg_reg[1]  (
	.SI(serialized_data),
	.SE(test_se),
	.RN(rst_n),
	.Q(parallel_data_reg[1]),
	.D(n33),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \parallel_data_reg_reg[7]  (
	.SI(parallel_data_reg[6]),
	.SE(test_se),
	.RN(rst_n),
	.Q(parallel_data_reg[7]),
	.D(n27),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \parallel_data_reg_reg[0]  (
	.SI(n35),
	.SE(test_se),
	.RN(rst_n),
	.Q(serialized_data),
	.D(n34),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \counter_reg[2]  (
	.SI(n36),
	.SE(test_se),
	.RN(rst_n),
	.QN(n12),
	.Q(n35),
	.D(N26),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(rst_n),
	.Q(\counter[0] ),
	.D(N24),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \counter_reg[1]  (
	.SI(\counter[0] ),
	.SE(test_se),
	.RN(rst_n),
	.QN(n13),
	.Q(n36),
	.D(N25),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U14 (
	.Y(n18),
	.B(n16),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U15 (
	.Y(n15),
	.B(n18),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U16 (
	.Y(n25),
	.B(serilaizer_enable),
	.AN(serilaizer_done), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U17 (
	.Y(n16),
	.B(busy),
	.AN(data_valid), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U18 (
	.Y(n34),
	.B0(n24),
	.A1N(n15),
	.A0N(serialized_data), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U19 (
	.Y(n24),
	.B1(n16),
	.B0(p_data[0]),
	.A1(n18),
	.A0(parallel_data_reg[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U20 (
	.Y(n33),
	.B0(n23),
	.A1N(parallel_data_reg[1]),
	.A0N(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U21 (
	.Y(n23),
	.B1(n16),
	.B0(p_data[1]),
	.A1(n18),
	.A0(parallel_data_reg[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U22 (
	.Y(n32),
	.B0(n22),
	.A1N(parallel_data_reg[2]),
	.A0N(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U23 (
	.Y(n22),
	.B1(n16),
	.B0(p_data[2]),
	.A1(n18),
	.A0(parallel_data_reg[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U24 (
	.Y(n31),
	.B0(n21),
	.A1N(parallel_data_reg[3]),
	.A0N(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U25 (
	.Y(n21),
	.B1(n16),
	.B0(p_data[3]),
	.A1(n18),
	.A0(parallel_data_reg[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U26 (
	.Y(n30),
	.B0(n20),
	.A1N(parallel_data_reg[4]),
	.A0N(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U27 (
	.Y(n20),
	.B1(n16),
	.B0(p_data[4]),
	.A1(n18),
	.A0(parallel_data_reg[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U28 (
	.Y(n29),
	.B0(n19),
	.A1N(parallel_data_reg[5]),
	.A0N(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U29 (
	.Y(n19),
	.B1(n16),
	.B0(p_data[5]),
	.A1(n18),
	.A0(parallel_data_reg[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U30 (
	.Y(n28),
	.B0(n17),
	.A1N(parallel_data_reg[6]),
	.A0N(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U31 (
	.Y(n17),
	.B1(n16),
	.B0(p_data[6]),
	.A1(parallel_data_reg[7]),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U32 (
	.Y(n27),
	.B1(n16),
	.B0(p_data[7]),
	.A1(parallel_data_reg[7]),
	.A0(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U33 (
	.Y(serilaizer_done),
	.C(n12),
	.B(n14),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U34 (
	.Y(N26),
	.B1(n25),
	.B0(n12),
	.A2(n13),
	.A1(n14),
	.A0(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U35 (
	.Y(N24),
	.B(n25),
	.A(\counter[0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U36 (
	.Y(N25),
	.B(n25),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U37 (
	.Y(n26),
	.B(\counter[0] ),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U38 (
	.Y(n14),
	.A(\counter[0] ), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module parity_calc_test_1 (
	p_data, 
	data_valid, 
	busy, 
	parity_type, 
	clk, 
	rst_n, 
	parity_bit, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input [7:0] p_data;
   input data_valid;
   input busy;
   input parity_type;
   input clk;
   input rst_n;
   output parity_bit;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n8;

   // Module instantiations
   SDFFRQX2M parity_bit_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(rst_n),
	.Q(parity_bit),
	.D(n8),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U2 (
	.Y(n5),
	.B(p_data[2]),
	.A(p_data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U3 (
	.Y(n3),
	.C(n6),
	.B(p_data[4]),
	.A(p_data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U4 (
	.Y(n6),
	.B(p_data[6]),
	.A(p_data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U5 (
	.Y(n8),
	.B1(n2),
	.B0(n1),
	.A1N(n2),
	.A0N(parity_bit), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U6 (
	.Y(n2),
	.B(data_valid),
	.AN(busy), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U7 (
	.Y(n1),
	.C(n4),
	.B(parity_type),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U8 (
	.Y(n4),
	.C(n5),
	.B(p_data[0]),
	.A(p_data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux (
	mux_sel, 
	parity_bit, 
	serialized_data, 
	tx_out, 
	VDD, 
	VSS);
   input [1:0] mux_sel;
   input parity_bit;
   input serialized_data;
   output tx_out;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n2;
   wire n1;
   wire n3;
   wire n4;
   wire n5;

   // Module instantiations
   AND3X2M U3 (
	.Y(n1),
	.C(serialized_data),
	.B(n5),
	.A(mux_sel[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX12M U4 (
	.Y(tx_out),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U5 (
	.Y(n4),
	.B(n5),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U6 (
	.Y(n3),
	.B(n1),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U7 (
	.Y(n5),
	.A(mux_sel[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U8 (
	.Y(n2),
	.B(parity_bit),
	.AN(mux_sel[1]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module rst_synchronizer_test_0 (
	clk, 
	rst_n, 
	sync_rst, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input clk;
   input rst_n;
   output sync_rst;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire [2:1] syn_rst_reg;

   assign test_so = syn_rst_reg[2] ;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \syn_rst_reg_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(rst_n),
	.Q(sync_rst),
	.D(syn_rst_reg[1]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \syn_rst_reg_reg[2]  (
	.SI(syn_rst_reg[1]),
	.SE(test_se),
	.RN(rst_n),
	.Q(syn_rst_reg[2]),
	.D(HTIE_LTIEHI_NET),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M \syn_rst_reg_reg[1]  (
	.SI(sync_rst),
	.SE(test_se),
	.RN(rst_n),
	.Q(syn_rst_reg[1]),
	.D(syn_rst_reg[2]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module rst_synchronizer_test_1 (
	clk, 
	rst_n, 
	sync_rst, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input clk;
   input rst_n;
   output sync_rst;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire [2:1] syn_rst_reg;

   assign test_so = syn_rst_reg[2] ;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \syn_rst_reg_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(rst_n),
	.Q(sync_rst),
	.D(syn_rst_reg[1]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \syn_rst_reg_reg[2]  (
	.SI(syn_rst_reg[1]),
	.SE(test_se),
	.RN(rst_n),
	.Q(syn_rst_reg[2]),
	.D(HTIE_LTIEHI_NET),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M \syn_rst_reg_reg[1]  (
	.SI(sync_rst),
	.SE(test_se),
	.RN(rst_n),
	.Q(syn_rst_reg[1]),
	.D(syn_rst_reg[2]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module clock_gating (
	clk_enable, 
	clk, 
	gated_clk, 
	VDD, 
	VSS);
   input clk_enable;
   input clk;
   output gated_clk;
   inout VDD;
   inout VSS;

   // Module instantiations
   TLATNCAX3M dut0 (
	.ECK(gated_clk),
	.E(clk_enable),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module clk_div_test_1 (
	i_ref_clk, 
	i_rst_n, 
	i_clk_en, 
	i_div_ratio, 
	o_div_clk, 
	test_si, 
	test_so, 
	test_se, 
	tx_clk__Exclude_0_NET, 
	scan_clk_uart_clk_mux_out__L6_N0, 
	scan_clk_uart_clk_mux_out__L6_N2, 
	VDD, 
	VSS);
   input i_ref_clk;
   input i_rst_n;
   input i_clk_en;
   input [7:0] i_div_ratio;
   output o_div_clk;
   input test_si;
   output test_so;
   input test_se;
   input tx_clk__Exclude_0_NET;
   input scan_clk_uart_clk_mux_out__L6_N0;
   input scan_clk_uart_clk_mux_out__L6_N2;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN8_n55;
   wire n16__Exclude_0_NET;
   wire HTIE_LTIEHI_NET;
   wire N8;
   wire N10;
   wire N11;
   wire N12;
   wire N13;
   wire N14;
   wire N15;
   wire N16;
   wire N17;
   wire n16;
   wire n19;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n17;
   wire n18;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire [7:0] counter;

   assign test_so = counter[7] ;

   // Module instantiations
   DLY3X1M FE_PHC8_n55 (
	.Y(n55),
	.A(FE_PHN8_n55), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX1M n16__Exclude_0 (
	.Y(n16__Exclude_0_NET),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M clk_reg_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(i_rst_n),
	.QN(n16),
	.Q(FE_PHN8_n55),
	.D(n25),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[4]  (
	.SI(counter[3]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[4]),
	.D(n30),
	.CK(scan_clk_uart_clk_mux_out__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[0]  (
	.SI(n55),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[0]),
	.D(n26),
	.CK(scan_clk_uart_clk_mux_out__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[6]  (
	.SI(counter[5]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[6]),
	.D(n32),
	.CK(scan_clk_uart_clk_mux_out__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[2]  (
	.SI(counter[1]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[2]),
	.D(n28),
	.CK(scan_clk_uart_clk_mux_out__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[5]  (
	.SI(counter[4]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[5]),
	.D(n31),
	.CK(scan_clk_uart_clk_mux_out__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[1]  (
	.SI(counter[0]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[1]),
	.D(n27),
	.CK(scan_clk_uart_clk_mux_out__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[3]  (
	.SI(counter[2]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[3]),
	.D(n29),
	.CK(scan_clk_uart_clk_mux_out__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[7]  (
	.SI(counter[6]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[7]),
	.D(n33),
	.CK(scan_clk_uart_clk_mux_out__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U19 (
	.Y(o_div_clk),
	.B1(n16),
	.B0(n19),
	.A1N(n19),
	.A0N(scan_clk_uart_clk_mux_out__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U4 (
	.Y(n1),
	.B(N8),
	.A(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U5 (
	.Y(n2),
	.B(N8),
	.A(counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U14 (
	.Y(n3),
	.B(N8),
	.A(counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U15 (
	.Y(n4),
	.B(N8),
	.A(counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U16 (
	.Y(n5),
	.B(N8),
	.A(counter[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U17 (
	.Y(n6),
	.B(N8),
	.A(counter[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U18 (
	.Y(n17),
	.B(N8),
	.A(counter[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U20 (
	.Y(n18),
	.B(counter[7]),
	.A(N8), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U21 (
	.Y(n19),
	.B(HTIE_LTIEHI_NET),
	.AN(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U22 (
	.Y(N8),
	.B(n46),
	.A(n45), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U23 (
	.Y(n33),
	.S0(n19),
	.B(counter[7]),
	.A(N17), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U24 (
	.Y(n32),
	.S0(n19),
	.B(counter[6]),
	.A(N16), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U25 (
	.Y(n31),
	.S0(n19),
	.B(counter[5]),
	.A(N15), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U26 (
	.Y(n30),
	.S0(n19),
	.B(counter[4]),
	.A(N14), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U27 (
	.Y(n29),
	.S0(n19),
	.B(counter[3]),
	.A(N13), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U28 (
	.Y(n28),
	.S0(n19),
	.B(counter[2]),
	.A(N12), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U29 (
	.Y(n27),
	.S0(n19),
	.B(counter[1]),
	.A(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U30 (
	.Y(n26),
	.S0(n19),
	.B(counter[0]),
	.A(N10), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U31 (
	.Y(n25),
	.S0(n19),
	.B(n16__Exclude_0_NET),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U32 (
	.Y(n20),
	.B(n21),
	.A(tx_clk__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U33 (
	.Y(n21),
	.C0(n35),
	.B1(n34),
	.B0(n24),
	.A1(n23),
	.A0(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U34 (
	.Y(n35),
	.A(N8), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U35 (
	.Y(n34),
	.D(n38),
	.C(n37),
	.B(n36),
	.A(counter[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U36 (
	.Y(n38),
	.B(counter[2]),
	.A(i_div_ratio[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U37 (
	.Y(n37),
	.B(counter[1]),
	.A(i_div_ratio[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U38 (
	.Y(n36),
	.B(counter[0]),
	.A(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U39 (
	.Y(n24),
	.D(n42),
	.C(n41),
	.B(n40),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U40 (
	.Y(n42),
	.B(counter[6]),
	.A(i_div_ratio[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U41 (
	.Y(n41),
	.B(counter[5]),
	.A(i_div_ratio[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U42 (
	.Y(n40),
	.B(counter[4]),
	.A(i_div_ratio[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U43 (
	.Y(n39),
	.B(counter[3]),
	.A(i_div_ratio[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U44 (
	.Y(n23),
	.D(counter[4]),
	.C(counter[5]),
	.B(counter[6]),
	.A(counter[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U45 (
	.Y(n22),
	.D(counter[0]),
	.C(counter[1]),
	.B(counter[2]),
	.A(counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4BX1M U46 (
	.Y(n43),
	.D(i_div_ratio[1]),
	.C(i_div_ratio[3]),
	.B(i_div_ratio[2]),
	.AN(n44), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U47 (
	.Y(n44),
	.D(i_div_ratio[4]),
	.C(i_div_ratio[5]),
	.B(i_div_ratio[6]),
	.A(i_div_ratio[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U48 (
	.Y(n46),
	.D(n50),
	.C(n49),
	.B(n48),
	.A(n47), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U49 (
	.Y(n50),
	.B(counter[7]),
	.A(i_div_ratio[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U50 (
	.Y(n49),
	.B(counter[2]),
	.A(i_div_ratio[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U51 (
	.Y(n48),
	.B(counter[1]),
	.A(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U52 (
	.Y(n47),
	.B(counter[0]),
	.A(i_div_ratio[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U53 (
	.Y(n45),
	.D(n54),
	.C(n53),
	.B(n52),
	.A(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U54 (
	.Y(n54),
	.B(counter[6]),
	.A(i_div_ratio[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U55 (
	.Y(n53),
	.B(counter[5]),
	.A(i_div_ratio[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U56 (
	.Y(n52),
	.B(counter[4]),
	.A(i_div_ratio[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U57 (
	.Y(n51),
	.B(counter[3]),
	.A(i_div_ratio[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   clk_div_0_DW01_inc_0 add_21_aco (
	.A({ n18,
		n17,
		n6,
		n5,
		n4,
		n3,
		n2,
		n1 }),
	.SUM({ N17,
		N16,
		N15,
		N14,
		N13,
		N12,
		N11,
		N10 }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module clk_div_0_DW01_inc_0 (
	A, 
	SUM, 
	VDD, 
	VSS);
   input [7:0] A;
   output [7:0] SUM;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [7:2] carry;

   // Module instantiations
   ADDHX1M U1_1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.B(carry[6]),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.B(carry[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.B(carry[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.B(carry[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.B(carry[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.B(A[0]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U1 (
	.Y(SUM[7]),
	.B(A[7]),
	.A(carry[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U2 (
	.Y(SUM[0]),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module clk_div_test_0 (
	i_ref_clk, 
	i_rst_n, 
	i_clk_en, 
	i_div_ratio, 
	o_div_clk, 
	test_si, 
	test_so, 
	test_se, 
	rx_clk__Exclude_0_NET, 
	scan_clk_uart_clk_mux_out__L6_N1, 
	scan_clk_uart_clk_mux_out__L6_N3, 
	VDD, 
	VSS);
   input i_ref_clk;
   input i_rst_n;
   input i_clk_en;
   input [7:0] i_div_ratio;
   output o_div_clk;
   input test_si;
   output test_so;
   input test_se;
   input rx_clk__Exclude_0_NET;
   input scan_clk_uart_clk_mux_out__L6_N1;
   input scan_clk_uart_clk_mux_out__L6_N3;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN7_n75;
   wire n65__Exclude_0_NET;
   wire HTIE_LTIEHI_NET;
   wire LTIE_LTIELO_NET;
   wire N8;
   wire N10;
   wire N11;
   wire N12;
   wire N13;
   wire N14;
   wire N15;
   wire N16;
   wire N17;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n17;
   wire n18;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n75;
   wire [7:0] counter;

   assign test_so = counter[7] ;

   // Module instantiations
   DLY2X1M FE_PHC7_n75 (
	.Y(n75),
	.A(FE_PHN7_n75), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX1M n65__Exclude_0 (
	.Y(n65__Exclude_0_NET),
	.A(n65), 
	.VDD(VDD), 
	.VSS(VSS));
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   TIELOM LTIE_LTIELO (
	.Y(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M clk_reg_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(i_rst_n),
	.QN(n65),
	.Q(FE_PHN7_n75),
	.D(n63),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[4]  (
	.SI(counter[3]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[4]),
	.D(n58),
	.CK(scan_clk_uart_clk_mux_out__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[0]  (
	.SI(n75),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[0]),
	.D(n62),
	.CK(scan_clk_uart_clk_mux_out__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[6]  (
	.SI(counter[5]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[6]),
	.D(n56),
	.CK(scan_clk_uart_clk_mux_out__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[2]  (
	.SI(counter[1]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[2]),
	.D(n60),
	.CK(scan_clk_uart_clk_mux_out__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[5]  (
	.SI(counter[4]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[5]),
	.D(n57),
	.CK(scan_clk_uart_clk_mux_out__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[1]  (
	.SI(counter[0]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[1]),
	.D(n61),
	.CK(scan_clk_uart_clk_mux_out__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[3]  (
	.SI(counter[2]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[3]),
	.D(n59),
	.CK(scan_clk_uart_clk_mux_out__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[7]  (
	.SI(counter[6]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[7]),
	.D(n55),
	.CK(scan_clk_uart_clk_mux_out__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U19 (
	.Y(o_div_clk),
	.B1(n65),
	.B0(n64),
	.A1N(n64),
	.A0N(scan_clk_uart_clk_mux_out__L6_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U4 (
	.Y(n1),
	.B(N8),
	.A(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U5 (
	.Y(n2),
	.B(N8),
	.A(counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U14 (
	.Y(n3),
	.B(N8),
	.A(counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U15 (
	.Y(n4),
	.B(N8),
	.A(counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U16 (
	.Y(n5),
	.B(N8),
	.A(counter[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U17 (
	.Y(n6),
	.B(N8),
	.A(counter[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U18 (
	.Y(n17),
	.B(N8),
	.A(counter[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U20 (
	.Y(n18),
	.B(counter[7]),
	.A(N8), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U21 (
	.Y(n64),
	.B(HTIE_LTIEHI_NET),
	.AN(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U22 (
	.Y(N8),
	.B(n46),
	.A(n45), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U23 (
	.Y(n55),
	.S0(n64),
	.B(counter[7]),
	.A(N17), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U24 (
	.Y(n56),
	.S0(n64),
	.B(counter[6]),
	.A(N16), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U25 (
	.Y(n57),
	.S0(n64),
	.B(counter[5]),
	.A(N15), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U26 (
	.Y(n58),
	.S0(n64),
	.B(counter[4]),
	.A(N14), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U27 (
	.Y(n59),
	.S0(n64),
	.B(counter[3]),
	.A(N13), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U28 (
	.Y(n60),
	.S0(n64),
	.B(counter[2]),
	.A(N12), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U29 (
	.Y(n61),
	.S0(n64),
	.B(counter[1]),
	.A(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U30 (
	.Y(n62),
	.S0(n64),
	.B(counter[0]),
	.A(N10), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U31 (
	.Y(n63),
	.S0(n64),
	.B(n65__Exclude_0_NET),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U32 (
	.Y(n20),
	.B(n21),
	.A(rx_clk__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U33 (
	.Y(n21),
	.C0(n35),
	.B1(n34),
	.B0(n24),
	.A1(n23),
	.A0(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U34 (
	.Y(n35),
	.A(N8), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U35 (
	.Y(n34),
	.D(n38),
	.C(n37),
	.B(n36),
	.A(counter[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U36 (
	.Y(n38),
	.B(counter[2]),
	.A(i_div_ratio[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U37 (
	.Y(n37),
	.B(counter[1]),
	.A(i_div_ratio[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U38 (
	.Y(n36),
	.B(counter[0]),
	.A(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U39 (
	.Y(n24),
	.D(n42),
	.C(n41),
	.B(n40),
	.A(n39), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U40 (
	.Y(n42),
	.B(counter[6]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U41 (
	.Y(n41),
	.B(counter[5]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U42 (
	.Y(n40),
	.B(counter[4]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U43 (
	.Y(n39),
	.B(counter[3]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U44 (
	.Y(n23),
	.D(counter[4]),
	.C(counter[5]),
	.B(counter[6]),
	.A(counter[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U45 (
	.Y(n22),
	.D(counter[0]),
	.C(counter[1]),
	.B(counter[2]),
	.A(counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4BX1M U46 (
	.Y(n43),
	.D(i_div_ratio[1]),
	.C(i_div_ratio[3]),
	.B(i_div_ratio[2]),
	.AN(n44), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U47 (
	.Y(n44),
	.D(LTIE_LTIELO_NET),
	.C(LTIE_LTIELO_NET),
	.B(LTIE_LTIELO_NET),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U48 (
	.Y(n46),
	.D(n50),
	.C(n49),
	.B(n48),
	.A(n47), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U49 (
	.Y(n50),
	.B(counter[7]),
	.A(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U50 (
	.Y(n49),
	.B(counter[2]),
	.A(i_div_ratio[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U51 (
	.Y(n48),
	.B(counter[1]),
	.A(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U52 (
	.Y(n47),
	.B(counter[0]),
	.A(i_div_ratio[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U53 (
	.Y(n45),
	.D(n42),
	.C(n41),
	.B(n40),
	.A(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U57 (
	.Y(n51),
	.B(counter[3]),
	.A(i_div_ratio[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   clk_div_1_DW01_inc_0 add_21_aco (
	.A({ n18,
		n17,
		n6,
		n5,
		n4,
		n3,
		n2,
		n1 }),
	.SUM({ N17,
		N16,
		N15,
		N14,
		N13,
		N12,
		N11,
		N10 }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module clk_div_1_DW01_inc_0 (
	A, 
	SUM, 
	VDD, 
	VSS);
   input [7:0] A;
   output [7:0] SUM;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [7:2] carry;

   // Module instantiations
   ADDHX1M U1_1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.B(carry[6]),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.B(carry[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.B(carry[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.B(carry[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.B(carry[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.B(A[0]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U1 (
	.Y(SUM[7]),
	.B(A[7]),
	.A(carry[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U2 (
	.Y(SUM[0]),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module pulse_gen_test_1 (
	clk, 
	rst_n, 
	in, 
	d2, 
	out, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input clk;
   input rst_n;
   input in;
   output d2;
   output out;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire q;

   assign test_so = q ;

   // Module instantiations
   SDFFRQX2M q_reg (
	.SI(out),
	.SE(test_se),
	.RN(rst_n),
	.Q(q),
	.D(in),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M out_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(rst_n),
	.Q(out),
	.D(d2),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U5 (
	.Y(d2),
	.B(q),
	.AN(in), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module system_TOP (
	Ref_clk, 
	Uart_clk, 
	rst_n, 
	rx_in, 
	tx_out, 
	stop_error, 
	parity_error, 
	start_glitch, 
	SI, 
	SE, 
	TESTMODE, 
	SCAN_CLK, 
	SCAN_RST, 
	SO, 
	VDD, 
	VSS);
   input Ref_clk;
   input Uart_clk;
   input rst_n;
   input rx_in;
   output tx_out;
   output stop_error;
   output parity_error;
   output start_glitch;
   input [4:0] SI;
   input SE;
   input TESTMODE;
   input SCAN_CLK;
   input SCAN_RST;
   output [4:0] SO;
   inout VDD;
   inout VSS;

   // Internal wires
   wire Ref_clk__L2_N0;
   wire Ref_clk__L1_N0;
   wire Uart_clk__L2_N0;
   wire Uart_clk__L1_N0;
   wire SCAN_CLK__L7_N0;
   wire SCAN_CLK__L6_N0;
   wire SCAN_CLK__L5_N1;
   wire SCAN_CLK__L5_N0;
   wire SCAN_CLK__L4_N0;
   wire SCAN_CLK__L3_N0;
   wire SCAN_CLK__L2_N1;
   wire SCAN_CLK__L2_N0;
   wire SCAN_CLK__L1_N0;
   wire scan_clk_uart_clk_mux_out__L6_N3;
   wire scan_clk_uart_clk_mux_out__L6_N2;
   wire scan_clk_uart_clk_mux_out__L6_N1;
   wire scan_clk_uart_clk_mux_out__L6_N0;
   wire scan_clk_uart_clk_mux_out__L5_N1;
   wire scan_clk_uart_clk_mux_out__L5_N0;
   wire scan_clk_uart_clk_mux_out__L4_N1;
   wire scan_clk_uart_clk_mux_out__L4_N0;
   wire scan_clk_uart_clk_mux_out__L3_N1;
   wire scan_clk_uart_clk_mux_out__L3_N0;
   wire scan_clk_uart_clk_mux_out__L2_N3;
   wire scan_clk_uart_clk_mux_out__L2_N2;
   wire scan_clk_uart_clk_mux_out__L2_N1;
   wire scan_clk_uart_clk_mux_out__L2_N0;
   wire scan_clk_uart_clk_mux_out__L1_N1;
   wire scan_clk_uart_clk_mux_out__L1_N0;
   wire tx_clk__Exclude_0_NET;
   wire rx_clk__Exclude_0_NET;
   wire scan_clk_ref_clk_mux_out__L4_N1;
   wire scan_clk_ref_clk_mux_out__L4_N0;
   wire scan_clk_ref_clk_mux_out__L3_N0;
   wire scan_clk_ref_clk_mux_out__L2_N0;
   wire scan_clk_ref_clk_mux_out__L1_N0;
   wire gated_clk__L1_N0;
   wire scan_clk_uart_tx_clk_mux_out__L1_N0;
   wire scan_clk_uart_rx_clk_mux_out__L1_N0;
   wire FE_OFN13_SE;
   wire FE_OFN6_scan_rst_sync2_mux_out;
   wire FE_OFN4_scan_rst_sync1_mux_out;
   wire FE_OFN3_scan_rst_sync1_mux_out;
   wire FE_OFN2_scan_rst_sync1_mux_out;
   wire FE_OFN0_scan_rst_sync1_mux_out;
   wire scan_clk_uart_clk_mux_out;
   wire scan_clk_ref_clk_mux_out;
   wire tx_clk;
   wire scan_clk_uart_tx_clk_mux_out;
   wire rx_clk;
   wire scan_clk_uart_rx_clk_mux_out;
   wire scan_rst_mux_out;
   wire ref_sync_rst;
   wire scan_rst_sync1_mux_out;
   wire uart_sync_rst;
   wire scan_rst_sync2_mux_out;
   wire empty_flag;
   wire q1;
   wire out_valid;
   wire rx_d_valid;
   wire full_flag;
   wire rd_data_valid;
   wire alu_en;
   wire clk_en;
   wire w_en;
   wire r_en;
   wire w_inc;
   wire data_valid;
   wire gated_clk;
   wire rd_inc;
   wire busy;
   wire _1_net_;
   wire n3;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n14;
   wire n15;
   wire n16;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n42;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire [7:0] reg2;
   wire [3:0] out;
   wire [15:0] alu_out;
   wire [7:0] rx_P_data;
   wire [7:0] rd_data;
   wire [3:0] alu_fun;
   wire [3:0] address;
   wire [7:0] w_data;
   wire [7:0] tx_P_data;
   wire [7:0] p_data;
   wire [7:0] reg0;
   wire [7:0] reg1;
   wire [7:0] reg3;
   wire [7:0] fifo_rd_data;

   assign SO[2] = reg2[3] ;

   // Module instantiations
   CLKINVX40M Ref_clk__L2_I0 (
	.Y(Ref_clk__L2_N0),
	.A(Ref_clk__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M Ref_clk__L1_I0 (
	.Y(Ref_clk__L1_N0),
	.A(Ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M Uart_clk__L2_I0 (
	.Y(Uart_clk__L2_N0),
	.A(Uart_clk__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M Uart_clk__L1_I0 (
	.Y(Uart_clk__L1_N0),
	.A(Uart_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M SCAN_CLK__L7_I0 (
	.Y(SCAN_CLK__L7_N0),
	.A(SCAN_CLK__L6_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX1M SCAN_CLK__L6_I0 (
	.Y(SCAN_CLK__L6_N0),
	.A(SCAN_CLK__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX5M SCAN_CLK__L5_I1 (
	.Y(SCAN_CLK__L5_N1),
	.A(SCAN_CLK__L4_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M SCAN_CLK__L5_I0 (
	.Y(SCAN_CLK__L5_N0),
	.A(SCAN_CLK__L4_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM SCAN_CLK__L4_I0 (
	.Y(SCAN_CLK__L4_N0),
	.A(SCAN_CLK__L3_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM SCAN_CLK__L3_I0 (
	.Y(SCAN_CLK__L3_N0),
	.A(SCAN_CLK__L2_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX1M SCAN_CLK__L2_I1 (
	.Y(SCAN_CLK__L2_N1),
	.A(SCAN_CLK__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M SCAN_CLK__L2_I0 (
	.Y(SCAN_CLK__L2_N0),
	.A(SCAN_CLK__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M SCAN_CLK__L1_I0 (
	.Y(SCAN_CLK__L1_N0),
	.A(SCAN_CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M scan_clk_uart_clk_mux_out__L6_I3 (
	.Y(scan_clk_uart_clk_mux_out__L6_N3),
	.A(scan_clk_uart_clk_mux_out__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M scan_clk_uart_clk_mux_out__L6_I2 (
	.Y(scan_clk_uart_clk_mux_out__L6_N2),
	.A(scan_clk_uart_clk_mux_out__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M scan_clk_uart_clk_mux_out__L6_I1 (
	.Y(scan_clk_uart_clk_mux_out__L6_N1),
	.A(scan_clk_uart_clk_mux_out__L5_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M scan_clk_uart_clk_mux_out__L6_I0 (
	.Y(scan_clk_uart_clk_mux_out__L6_N0),
	.A(scan_clk_uart_clk_mux_out__L5_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M scan_clk_uart_clk_mux_out__L5_I1 (
	.Y(scan_clk_uart_clk_mux_out__L5_N1),
	.A(scan_clk_uart_clk_mux_out__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M scan_clk_uart_clk_mux_out__L5_I0 (
	.Y(scan_clk_uart_clk_mux_out__L5_N0),
	.A(scan_clk_uart_clk_mux_out__L4_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M scan_clk_uart_clk_mux_out__L4_I1 (
	.Y(scan_clk_uart_clk_mux_out__L4_N1),
	.A(scan_clk_uart_clk_mux_out__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M scan_clk_uart_clk_mux_out__L4_I0 (
	.Y(scan_clk_uart_clk_mux_out__L4_N0),
	.A(scan_clk_uart_clk_mux_out__L3_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM scan_clk_uart_clk_mux_out__L3_I1 (
	.Y(scan_clk_uart_clk_mux_out__L3_N1),
	.A(scan_clk_uart_clk_mux_out__L2_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M scan_clk_uart_clk_mux_out__L3_I0 (
	.Y(scan_clk_uart_clk_mux_out__L3_N0),
	.A(scan_clk_uart_clk_mux_out__L2_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM scan_clk_uart_clk_mux_out__L2_I3 (
	.Y(scan_clk_uart_clk_mux_out__L2_N3),
	.A(scan_clk_uart_clk_mux_out__L1_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M scan_clk_uart_clk_mux_out__L2_I2 (
	.Y(scan_clk_uart_clk_mux_out__L2_N2),
	.A(scan_clk_uart_clk_mux_out__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M scan_clk_uart_clk_mux_out__L2_I1 (
	.Y(scan_clk_uart_clk_mux_out__L2_N1),
	.A(scan_clk_uart_clk_mux_out__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX4M scan_clk_uart_clk_mux_out__L2_I0 (
	.Y(scan_clk_uart_clk_mux_out__L2_N0),
	.A(scan_clk_uart_clk_mux_out__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M scan_clk_uart_clk_mux_out__L1_I1 (
	.Y(scan_clk_uart_clk_mux_out__L1_N1),
	.A(scan_clk_uart_clk_mux_out), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX32M scan_clk_uart_clk_mux_out__L1_I0 (
	.Y(scan_clk_uart_clk_mux_out__L1_N0),
	.A(scan_clk_uart_clk_mux_out), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX1M tx_clk__Exclude_0 (
	.Y(tx_clk__Exclude_0_NET),
	.A(tx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX1M rx_clk__Exclude_0 (
	.Y(rx_clk__Exclude_0_NET),
	.A(rx_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M scan_clk_ref_clk_mux_out__L4_I1 (
	.Y(scan_clk_ref_clk_mux_out__L4_N1),
	.A(scan_clk_ref_clk_mux_out__L3_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M scan_clk_ref_clk_mux_out__L4_I0 (
	.Y(scan_clk_ref_clk_mux_out__L4_N0),
	.A(scan_clk_ref_clk_mux_out__L3_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX40M scan_clk_ref_clk_mux_out__L3_I0 (
	.Y(scan_clk_ref_clk_mux_out__L3_N0),
	.A(scan_clk_ref_clk_mux_out__L2_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M scan_clk_ref_clk_mux_out__L2_I0 (
	.Y(scan_clk_ref_clk_mux_out__L2_N0),
	.A(scan_clk_ref_clk_mux_out__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M scan_clk_ref_clk_mux_out__L1_I0 (
	.Y(scan_clk_ref_clk_mux_out__L1_N0),
	.A(scan_clk_ref_clk_mux_out), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M gated_clk__L1_I0 (
	.Y(gated_clk__L1_N0),
	.A(gated_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX16M scan_clk_uart_tx_clk_mux_out__L1_I0 (
	.Y(scan_clk_uart_tx_clk_mux_out__L1_N0),
	.A(scan_clk_uart_tx_clk_mux_out), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M scan_clk_uart_rx_clk_mux_out__L1_I0 (
	.Y(scan_clk_uart_rx_clk_mux_out__L1_N0),
	.A(scan_clk_uart_rx_clk_mux_out), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX4M FE_OFC13_SE (
	.Y(FE_OFN13_SE),
	.A(SE), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX8M FE_OFC6_scan_rst_sync2_mux_out (
	.Y(FE_OFN6_scan_rst_sync2_mux_out),
	.A(scan_rst_sync2_mux_out), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX8M FE_OFC4_scan_rst_sync1_mux_out (
	.Y(FE_OFN4_scan_rst_sync1_mux_out),
	.A(FE_OFN0_scan_rst_sync1_mux_out), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX8M FE_OFC3_scan_rst_sync1_mux_out (
	.Y(FE_OFN3_scan_rst_sync1_mux_out),
	.A(FE_OFN0_scan_rst_sync1_mux_out), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX8M FE_OFC2_scan_rst_sync1_mux_out (
	.Y(FE_OFN2_scan_rst_sync1_mux_out),
	.A(FE_OFN0_scan_rst_sync1_mux_out), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M FE_OFC0_scan_rst_sync1_mux_out (
	.Y(FE_OFN0_scan_rst_sync1_mux_out),
	.A(scan_rst_sync1_mux_out), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M q1_reg (
	.SI(n36),
	.SE(n52),
	.RN(FE_OFN6_scan_rst_sync2_mux_out),
	.Q(q1),
	.D(empty_flag),
	.CK(scan_clk_uart_tx_clk_mux_out__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M q2_reg (
	.SI(q1),
	.SE(n56),
	.RN(FE_OFN6_scan_rst_sync2_mux_out),
	.QN(n3),
	.Q(n35),
	.D(q1),
	.CK(scan_clk_uart_tx_clk_mux_out__L1_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U21 (
	.Y(_1_net_),
	.B(clk_en),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U22 (
	.Y(n9),
	.D(n21),
	.C(n22),
	.B(reg2[5]),
	.AN(reg2[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U23 (
	.Y(n10),
	.D(n21),
	.C(n22),
	.B(reg2[6]),
	.AN(reg2[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U24 (
	.Y(out[2]),
	.C(reg2[2]),
	.B(n46),
	.A(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U25 (
	.Y(out[1]),
	.C(reg2[2]),
	.B(n46),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U26 (
	.Y(out[3]),
	.D(reg2[6]),
	.C(reg2[7]),
	.B(reg2[5]),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U27 (
	.Y(n8),
	.C(reg2[4]),
	.B(n23),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U28 (
	.Y(out[0]),
	.C0(n23),
	.B0(n24),
	.A1(n12),
	.A0(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U29 (
	.Y(n11),
	.D(n22),
	.C(reg2[5]),
	.B(reg2[6]),
	.A(reg2[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U30 (
	.Y(n12),
	.B(n9),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U31 (
	.Y(n22),
	.A(reg2[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U32 (
	.Y(n23),
	.A(n46), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U33 (
	.Y(n24),
	.A(reg2[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U34 (
	.Y(n21),
	.A(reg2[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX4M U35 (
	.Y(n16),
	.A(address[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX4M U36 (
	.Y(n15),
	.A(address[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M U40 (
	.Y(n14),
	.A(TESTMODE), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX40M U42 (
	.Y(stop_error),
	.A(SO[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U43 (
	.Y(n45),
	.A(reg2[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U44 (
	.Y(n46),
	.A(n45), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U45 (
	.Y(n47),
	.A(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U46 (
	.Y(n48),
	.A(n58), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U47 (
	.Y(n49),
	.A(n48), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U48 (
	.Y(n50),
	.A(n48), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U49 (
	.Y(n51),
	.A(n59), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U50 (
	.Y(n52),
	.A(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U51 (
	.Y(n53),
	.A(n49), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U52 (
	.Y(n54),
	.A(n53), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U53 (
	.Y(n55),
	.A(FE_OFN13_SE), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U54 (
	.Y(n56),
	.A(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U55 (
	.Y(n57),
	.A(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   INVXLM U56 (
	.Y(n58),
	.A(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U57 (
	.Y(n59),
	.A(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   mux_2x1_0 scan_clk_uart_clk_mux (
	.in0(Uart_clk__L2_N0),
	.in1(SCAN_CLK__L2_N0),
	.sel(n14),
	.out(scan_clk_uart_clk_mux_out), 
	.VDD(VDD), 
	.VSS(VSS));
   mux_2x1_6 scan_clk_ref_clk_mux (
	.in0(Ref_clk__L2_N0),
	.in1(SCAN_CLK__L5_N0),
	.sel(n14),
	.out(scan_clk_ref_clk_mux_out), 
	.VDD(VDD), 
	.VSS(VSS));
   mux_2x1_5 scan_clk_uart_tx_clk_mux (
	.in0(tx_clk),
	.in1(SCAN_CLK__L7_N0),
	.sel(n14),
	.out(scan_clk_uart_tx_clk_mux_out), 
	.VDD(VDD), 
	.VSS(VSS));
   mux_2x1_4 scan_clk_uart_rx_clk_mux (
	.in0(rx_clk),
	.in1(SCAN_CLK__L7_N0),
	.sel(n14),
	.out(scan_clk_uart_rx_clk_mux_out), 
	.VDD(VDD), 
	.VSS(VSS));
   mux_2x1_3 scan_rst_mux (
	.in0(rst_n),
	.in1(SCAN_RST),
	.sel(n14),
	.out(scan_rst_mux_out), 
	.VDD(VDD), 
	.VSS(VSS));
   mux_2x1_2 scan_rst1_mux (
	.in0(ref_sync_rst),
	.in1(SCAN_RST),
	.sel(n14),
	.out(scan_rst_sync1_mux_out), 
	.VDD(VDD), 
	.VSS(VSS));
   mux_2x1_1 scan_rst2_mux (
	.in0(uart_sync_rst),
	.in1(SCAN_RST),
	.sel(n14),
	.out(scan_rst_sync2_mux_out), 
	.VDD(VDD), 
	.VSS(VSS));
   sys_ctrl_test_1 sys_ctrl (
	.clk(scan_clk_ref_clk_mux_out__L4_N0),
	.rst_n(scan_rst_sync1_mux_out),
	.alu_out({ alu_out[15],
		alu_out[14],
		alu_out[13],
		alu_out[12],
		alu_out[11],
		alu_out[10],
		alu_out[9],
		alu_out[8],
		alu_out[7],
		alu_out[6],
		alu_out[5],
		alu_out[4],
		alu_out[3],
		alu_out[2],
		alu_out[1],
		alu_out[0] }),
	.out_valid(out_valid),
	.rx_P_data({ rx_P_data[7],
		rx_P_data[6],
		rx_P_data[5],
		rx_P_data[4],
		rx_P_data[3],
		rx_P_data[2],
		rx_P_data[1],
		rx_P_data[0] }),
	.rx_d_valid(rx_d_valid),
	.full_flag(full_flag),
	.rd_data({ rd_data[7],
		rd_data[6],
		rd_data[5],
		rd_data[4],
		rd_data[3],
		rd_data[2],
		rd_data[1],
		rd_data[0] }),
	.rd_data_valid(rd_data_valid),
	.alu_en(alu_en),
	.alu_fun({ alu_fun[3],
		alu_fun[2],
		alu_fun[1],
		alu_fun[0] }),
	.clk_en(clk_en),
	.address({ address[3],
		address[2],
		address[1],
		address[0] }),
	.w_en(w_en),
	.r_en(r_en),
	.w_data({ w_data[7],
		w_data[6],
		w_data[5],
		w_data[4],
		w_data[3],
		w_data[2],
		w_data[1],
		w_data[0] }),
	.tx_P_data({ tx_P_data[7],
		tx_P_data[6],
		tx_P_data[5],
		tx_P_data[4],
		tx_P_data[3],
		tx_P_data[2],
		tx_P_data[1],
		tx_P_data[0] }),
	.w_inc(w_inc),
	.test_si(n29),
	.test_so(n28),
	.test_se(n57),
	.FE_OFN2_scan_rst_sync1_mux_out(FE_OFN2_scan_rst_sync1_mux_out), 
	.VDD(VDD), 
	.VSS(VSS));
   data_sync_top_module_test_1 data_sync (
	.dest_clk(scan_clk_ref_clk_mux_out__L4_N0),
	.dest_rst_n(FE_OFN2_scan_rst_sync1_mux_out),
	.unsync_bus({ p_data[7],
		p_data[6],
		p_data[5],
		p_data[4],
		p_data[3],
		p_data[2],
		p_data[1],
		p_data[0] }),
	.bus_enable(data_valid),
	.sync_bus({ rx_P_data[7],
		rx_P_data[6],
		rx_P_data[5],
		rx_P_data[4],
		rx_P_data[3],
		rx_P_data[2],
		rx_P_data[1],
		rx_P_data[0] }),
	.enable_pulse(rx_d_valid),
	.test_si(n37),
	.test_se(n52), 
	.VDD(VDD), 
	.VSS(VSS));
   RX_TOP_MODULE_test_1 uart_RX (
	.rx_in(rx_in),
	.prescale({ reg2[7],
		reg2[6],
		reg2[5],
		reg2[4],
		n46,
		reg2[2] }),
	.parity_enable(reg2[0]),
	.parity_type(reg2[1]),
	.rx_clk(scan_clk_uart_rx_clk_mux_out__L1_N0),
	.rst_n(FE_OFN6_scan_rst_sync2_mux_out),
	.p_data({ p_data[7],
		p_data[6],
		p_data[5],
		p_data[4],
		p_data[3],
		p_data[2],
		p_data[1],
		p_data[0] }),
	.stop_error(SO[0]),
	.parity_error(parity_error),
	.start_glitch(start_glitch),
	.data_valid(data_valid),
	.test_si2(n26),
	.test_si1(n27),
	.test_se(n47),
	.n23(n23),
	.FE_PT1_n24(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   RF_test_1 register_file (
	.wren(w_en),
	.rden(r_en),
	.clk(scan_clk_ref_clk_mux_out__L4_N0),
	.rst(scan_rst_sync1_mux_out),
	.wrdata({ w_data[7],
		w_data[6],
		w_data[5],
		w_data[4],
		w_data[3],
		w_data[2],
		w_data[1],
		w_data[0] }),
	.address({ address[3],
		address[2],
		n16,
		n15 }),
	.rddata({ rd_data[7],
		rd_data[6],
		rd_data[5],
		rd_data[4],
		rd_data[3],
		rd_data[2],
		rd_data[1],
		rd_data[0] }),
	.rddata_valid(rd_data_valid),
	.reg0({ reg0[7],
		reg0[6],
		reg0[5],
		reg0[4],
		reg0[3],
		reg0[2],
		reg0[1],
		reg0[0] }),
	.reg1({ reg1[7],
		reg1[6],
		reg1[5],
		reg1[4],
		reg1[3],
		reg1[2],
		reg1[1],
		reg1[0] }),
	.reg2({ reg2[7],
		reg2[6],
		reg2[5],
		reg2[4],
		reg2[3],
		reg2[2],
		reg2[1],
		reg2[0] }),
	.reg3({ reg3[7],
		reg3[6],
		reg3[5],
		reg3[4],
		reg3[3],
		reg3[2],
		reg3[1],
		reg3[0] }),
	.test_si3(SI[0]),
	.test_si2(SI[1]),
	.test_si1(n34),
	.test_so2(n30),
	.test_so1(SO[1]),
	.test_se(FE_OFN13_SE),
	.FE_OFN0_scan_rst_sync1_mux_out(FE_OFN0_scan_rst_sync1_mux_out),
	.FE_OFN2_scan_rst_sync1_mux_out(FE_OFN2_scan_rst_sync1_mux_out),
	.scan_clk_ref_clk_mux_out__L4_N1(scan_clk_ref_clk_mux_out__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   bit16_alu_test_1 alu (
	.a({ reg0[7],
		reg0[6],
		reg0[5],
		reg0[4],
		reg0[3],
		reg0[2],
		reg0[1],
		reg0[0] }),
	.b({ reg1[7],
		reg1[6],
		reg1[5],
		reg1[4],
		reg1[3],
		reg1[2],
		reg1[1],
		reg1[0] }),
	.alu_fun({ alu_fun[3],
		alu_fun[2],
		alu_fun[1],
		alu_fun[0] }),
	.clk(gated_clk__L1_N0),
	.rst_n(FE_OFN2_scan_rst_sync1_mux_out),
	.enable(alu_en),
	.alu_out({ alu_out[15],
		alu_out[14],
		alu_out[13],
		alu_out[12],
		alu_out[11],
		alu_out[10],
		alu_out[9],
		alu_out[8],
		alu_out[7],
		alu_out[6],
		alu_out[5],
		alu_out[4],
		alu_out[3],
		alu_out[2],
		alu_out[1],
		alu_out[0] }),
	.out_valid(out_valid),
	.test_si(n42),
	.test_se(n54),
	.FE_OFN3_scan_rst_sync1_mux_out(FE_OFN3_scan_rst_sync1_mux_out),
	.FE_OFN4_scan_rst_sync1_mux_out(FE_OFN4_scan_rst_sync1_mux_out), 
	.VDD(VDD), 
	.VSS(VSS));
   fifo_top_test_1 async_fifo (
	.w_clk(scan_clk_ref_clk_mux_out__L4_N0),
	.w_rst_n(FE_OFN2_scan_rst_sync1_mux_out),
	.rd_clk(scan_clk_uart_tx_clk_mux_out__L1_N0),
	.rd_rst_n(FE_OFN6_scan_rst_sync2_mux_out),
	.w_inc(w_inc),
	.rd_inc(rd_inc),
	.w_data({ tx_P_data[7],
		tx_P_data[6],
		tx_P_data[5],
		tx_P_data[4],
		tx_P_data[3],
		tx_P_data[2],
		tx_P_data[1],
		tx_P_data[0] }),
	.rd_data({ fifo_rd_data[7],
		fifo_rd_data[6],
		fifo_rd_data[5],
		fifo_rd_data[4],
		fifo_rd_data[3],
		fifo_rd_data[2],
		fifo_rd_data[1],
		fifo_rd_data[0] }),
	.full_flag(full_flag),
	.empty_flag(empty_flag),
	.test_si3(SI[2]),
	.test_si2(SI[3]),
	.test_si1(out_valid),
	.test_so3(n37),
	.test_so2(SO[3]),
	.test_so1(SO[4]),
	.test_se(FE_OFN13_SE),
	.FE_OFN3_scan_rst_sync1_mux_out(FE_OFN3_scan_rst_sync1_mux_out),
	.FE_OFN4_scan_rst_sync1_mux_out(FE_OFN4_scan_rst_sync1_mux_out),
	.scan_clk_ref_clk_mux_out__L4_N1(scan_clk_ref_clk_mux_out__L4_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   UART_tx_TOP_MODULE_test_1 UART_tx (
	.p_data({ fifo_rd_data[7],
		fifo_rd_data[6],
		fifo_rd_data[5],
		fifo_rd_data[4],
		fifo_rd_data[3],
		fifo_rd_data[2],
		fifo_rd_data[1],
		fifo_rd_data[0] }),
	.clk(scan_clk_uart_tx_clk_mux_out__L1_N0),
	.rst_n(FE_OFN6_scan_rst_sync2_mux_out),
	.data_valid(n3),
	.parity_type(reg2[1]),
	.parity_enable(reg2[0]),
	.tx_out(tx_out),
	.busy(busy),
	.test_si(SI[4]),
	.test_so(n42),
	.test_se(n56), 
	.VDD(VDD), 
	.VSS(VSS));
   rst_synchronizer_test_0 ref_clk_rst_sync (
	.clk(scan_clk_ref_clk_mux_out__L4_N0),
	.rst_n(scan_rst_mux_out),
	.sync_rst(ref_sync_rst),
	.test_si(n35),
	.test_so(n34),
	.test_se(n52), 
	.VDD(VDD), 
	.VSS(VSS));
   rst_synchronizer_test_1 uart_clk_rst_sync (
	.clk(scan_clk_uart_clk_mux_out__L6_N2),
	.rst_n(scan_rst_mux_out),
	.sync_rst(uart_sync_rst),
	.test_si(parity_error),
	.test_so(n26),
	.test_se(n59), 
	.VDD(VDD), 
	.VSS(VSS));
   clock_gating clock_gating_cell (
	.clk_enable(_1_net_),
	.clk(scan_clk_ref_clk_mux_out),
	.gated_clk(gated_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   clk_div_test_1 tx_div (
	.i_ref_clk(scan_clk_uart_clk_mux_out__L2_N0),
	.i_rst_n(scan_rst_sync2_mux_out),
	.i_clk_en(1'b1),
	.i_div_ratio({ reg3[7],
		reg3[6],
		reg3[5],
		reg3[4],
		reg3[3],
		reg3[2],
		reg3[1],
		reg3[0] }),
	.o_div_clk(tx_clk),
	.test_si(n28),
	.test_so(n27),
	.test_se(n59),
	.tx_clk__Exclude_0_NET(tx_clk__Exclude_0_NET),
	.scan_clk_uart_clk_mux_out__L6_N0(scan_clk_uart_clk_mux_out__L6_N0),
	.scan_clk_uart_clk_mux_out__L6_N2(scan_clk_uart_clk_mux_out__L6_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   clk_div_test_0 rx_div (
	.i_ref_clk(scan_clk_uart_clk_mux_out__L2_N1),
	.i_rst_n(scan_rst_sync2_mux_out),
	.i_clk_en(1'b1),
	.i_div_ratio({ 1'b0,
		1'b0,
		1'b0,
		1'b0,
		out[3],
		out[2],
		out[1],
		out[0] }),
	.o_div_clk(rx_clk),
	.test_si(n30),
	.test_so(n29),
	.test_se(n49),
	.rx_clk__Exclude_0_NET(rx_clk__Exclude_0_NET),
	.scan_clk_uart_clk_mux_out__L6_N1(scan_clk_uart_clk_mux_out__L6_N1),
	.scan_clk_uart_clk_mux_out__L6_N3(scan_clk_uart_clk_mux_out__L6_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   pulse_gen_test_1 pulse_gen (
	.clk(scan_clk_uart_tx_clk_mux_out__L1_N0),
	.rst_n(FE_OFN6_scan_rst_sync2_mux_out),
	.in(busy),
	.d2(rd_inc),
	.test_si(rx_P_data[7]),
	.test_so(n36),
	.test_se(n57), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

