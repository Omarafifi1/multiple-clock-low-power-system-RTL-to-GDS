

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO SYS_TOP 
  PIN SI[3] 
    ANTENNAPARTIALMETALAREA 0.269 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.29389 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.862 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.14862 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 18.344 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 88.427 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 461.313 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 2229.89 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.70919 LAYER VIA56 ;
  END SI[3]
  PIN SI[2] 
    ANTENNAPARTIALMETALAREA 0.629 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.02549 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.452 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.17652 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 2.6 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.6984 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 60.2251 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 297.046 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.03189 LAYER VIA45 ;
  END SI[2]
  PIN SI[1] 
    ANTENNAPARTIALMETALAREA 0.415 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.99615 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 3.256 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.8538 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 17.032 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 82.1163 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNAPARTIALMETALAREA 7.602 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 36.758 LAYER METAL6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL6 ; 
    ANTENNAMAXAREACAR 274.615 LAYER METAL6 ;
    ANTENNAMAXSIDEAREACAR 1335.48 LAYER METAL6 ;
    ANTENNAMAXCUTCAR 3.38649 LAYER VIA67 ;
  END SI[1]
  PIN SI[0] 
    ANTENNAPARTIALMETALAREA 1.028 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 5.13708 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 27.938 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 134.574 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 1.288 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.38768 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNAPARTIALMETALAREA 17.196 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 82.9052 LAYER METAL6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL6 ; 
    ANTENNAMAXAREACAR 336.529 LAYER METAL6 ;
    ANTENNAMAXSIDEAREACAR 1633.29 LAYER METAL6 ;
    ANTENNAMAXCUTCAR 3.38649 LAYER VIA67 ;
  END SI[0]
  PIN SO[3] 
    ANTENNAPARTIALMETALAREA 0.199 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.95719 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 17.278 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 83.2996 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNAPARTIALMETALAREA 7.5378 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 36.2241 LAYER METAL6 ;
    ANTENNAPARTIALCUTAREA 0.1296 LAYER VIA67 ;
    ANTENNADIFFAREA 0.537 LAYER METAL7 ; 
    ANTENNAPARTIALMETALAREA 40.74 LAYER METAL7 ;
    ANTENNAPARTIALMETALSIDEAREA 239.265 LAYER METAL7 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.221 LAYER METAL7 ; 
    ANTENNAMAXAREACAR 275.359 LAYER METAL7 ;
    ANTENNAMAXSIDEAREACAR 1531.59 LAYER METAL7 ;
  END SO[3]
  PIN SO[2] 
    ANTENNADIFFAREA 0.333 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 5.606 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.9649 LAYER METAL3 ;
  END SO[2]
  PIN SO[1] 
    ANTENNADIFFAREA 4.19 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 2.572 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.3713 LAYER METAL3 ;
  END SO[1]
  PIN SO[0] 
    ANTENNAPARTIALMETALAREA 41.252 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 198.615 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 3.748 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 18.2203 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.333 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 0.386 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.04906 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2002 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 78.3886 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 379.346 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.721279 LAYER VIA56 ;
  END SO[0]
  PIN scan_clk 
    ANTENNAPARTIALMETALAREA 0.255 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.22655 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 7.602 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 36.758 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 1.37 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.7821 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 1.61865 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 7.93145 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.0353598 LAYER VIA45 ;
  END scan_clk
  PIN scan_rst 
    ANTENNAPARTIALMETALAREA 0.387 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.86147 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 3.256 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.8538 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 18.238 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 88.1096 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1066 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 201.895 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 976.673 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 2.03189 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 3.748 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 18.2203 LAYER METAL5 ;
    ANTENNAGATEAREA 0.1599 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 225.335 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 1090.62 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.70919 LAYER VIA56 ;
  END scan_rst
  PIN test_mode 
    ANTENNAPARTIALMETALAREA 0.287 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.38047 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.878 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.41558 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 1.124 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.59884 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNAPARTIALMETALAREA 8.176 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 39.519 LAYER METAL6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.9279 LAYER METAL6 ; 
    ANTENNAMAXAREACAR 47.9385 LAYER METAL6 ;
    ANTENNAMAXSIDEAREACAR 234.866 LAYER METAL6 ;
    ANTENNAMAXCUTCAR 1.22026 LAYER VIA67 ;
  END test_mode
  PIN SE 
    ANTENNAPARTIALMETALAREA 0.273 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.31313 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.288 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.38768 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1157 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 14.5225 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 72.6213 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.936041 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 6.059 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 29.9134 LAYER METAL4 ;
    ANTENNAGATEAREA 2.314 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 32.8185 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 159.96 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 1.07125 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 6.406 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 31.3901 LAYER METAL5 ;
    ANTENNAGATEAREA 3.2994 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 34.7601 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 169.474 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 1.24806 LAYER VIA56 ;
  END SE
  PIN RST_N 
    ANTENNAPARTIALMETALAREA 0.975 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 4.68975 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.272 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.1207 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 3.912 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 19.0091 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 5.2 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 25.3968 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 174.709 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 854.934 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.70919 LAYER VIA56 ;
  END RST_N
  PIN UART_CLK 
    ANTENNAPARTIALMETALAREA 0.351 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.68831 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.632 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 3.23232 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.796 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.02116 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 0.628053 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 3.16668 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.0353598 LAYER VIA45 ;
  END UART_CLK
  PIN REF_CLK 
    ANTENNAPARTIALMETALAREA 0.291 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.39971 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.96 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.81 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 0.895782 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 4.45446 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.0353598 LAYER VIA45 ;
  END REF_CLK
  PIN UART_RX_IN 
    ANTENNAPARTIALMETALAREA 0.207 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.99567 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.355 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.70995 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 3.42 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 16.6426 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 12.03 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 58.0567 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNAPARTIALMETALAREA 3.256 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 15.8538 LAYER METAL6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.4693 LAYER METAL6 ; 
    ANTENNAMAXAREACAR 47.3293 LAYER METAL6 ;
    ANTENNAMAXSIDEAREACAR 231.267 LAYER METAL6 ;
    ANTENNAMAXCUTCAR 1.83108 LAYER VIA67 ;
  END UART_RX_IN
  PIN UART_TX_O 
    ANTENNADIFFAREA 0.861 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 2.326 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.1881 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.9347 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 5.65615 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 26.4249 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.077244 LAYER VIA34 ;
  END UART_TX_O
  PIN parity_error 
    ANTENNAPARTIALMETALAREA 0.199 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.95719 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 6.561 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 31.7508 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.537 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 25.97 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 125.108 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2405 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 133.31 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 647.487 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.11124 LAYER VIA56 ;
  END parity_error
  PIN framing_error 
    ANTENNAPARTIALMETALAREA 3.435 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.5224 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 0.537 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 18.098 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 87.2438 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2405 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 151.556 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 738.232 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.88401 LAYER VIA56 ;
  END framing_error
END SYS_TOP

END LIBRARY
