

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO system_TOP 
  PIN SI[4] 
    ANTENNAPARTIALMETALAREA 1.881 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.04761 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.878 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 4.41558 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 4.158 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 20.1924 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 16.622 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 80.1442 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 431.682 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 2090.18 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.70919 LAYER VIA56 ;
  END SI[4]
  PIN SI[3] 
    ANTENNAPARTIALMETALAREA 2.013 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.68253 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 1.862 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.14862 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 27.036 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 130.236 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 645.528 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 3118.78 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.70919 LAYER VIA56 ;
  END SI[3]
  PIN SI[2] 
    ANTENNAPARTIALMETALAREA 5.377 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 26.2482 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 103.502 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 504.412 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.677298 LAYER VIA23 ;
  END SI[2]
  PIN SI[1] 
    ANTENNAPARTIALMETALAREA 0.775 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 3.72775 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 4.814 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 23.3477 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 3.912 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 19.0091 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 1.862 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 9.14862 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 145.528 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 713.778 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.70919 LAYER VIA56 ;
  END SI[1]
  PIN SI[0] 
    ANTENNAPARTIALMETALAREA 0.233 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.12073 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 10.144 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 48.985 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 10.284 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 49.8508 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 225.528 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 1098.58 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.03189 LAYER VIA45 ;
  END SI[0]
  PIN SO[4] 
    ANTENNADIFFAREA 1.737 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 8.838 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 42.8956 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0702 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 134.725 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 653.944 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 1.54274 LAYER VIA34 ;
  END SO[4]
  PIN SO[3] 
    ANTENNADIFFAREA 1.737 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 2.138 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.4762 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0702 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 72.4031 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 351.435 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 1.54274 LAYER VIA34 ;
  END SO[3]
  PIN SO[2] 
    ANTENNAPARTIALMETALAREA 0.194 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.93314 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 5.599 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 27.1236 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 1.737 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 32.202 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 155.084 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1404 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 329.405 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 1590.35 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.05698 LAYER VIA56 ;
  END SO[2]
  PIN SO[1] 
    ANTENNAPARTIALMETALAREA 0.199 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.95719 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 2.419 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.8278 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 25.806 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 124.319 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNADIFFAREA 1.737 LAYER METAL6 ; 
    ANTENNAPARTIALMETALAREA 9.956 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 48.2732 LAYER METAL6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0702 LAYER METAL6 ; 
    ANTENNAMAXAREACAR 175.195 LAYER METAL6 ;
    ANTENNAMAXSIDEAREACAR 859.569 LAYER METAL6 ;
    ANTENNAMAXCUTCAR 2.57123 LAYER VIA67 ;
  END SO[1]
  PIN SO[0] 
    ANTENNAPARTIALMETALAREA 37.978 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 182.867 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNADIFFAREA 1.431 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 25.372 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 122.424 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0192 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 64.5923 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 316.95 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 1.70888 LAYER VIA45 ;
  END SO[0]
  PIN Ref_clk 
    ANTENNAPARTIALMETALAREA 0.291 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.39971 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.222 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.26022 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 3.888 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 19.0861 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 1.85177 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 9.11558 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.0353598 LAYER VIA45 ;
  END Ref_clk
  PIN Uart_clk 
    ANTENNAPARTIALMETALAREA 0.269 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.29389 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 18.098 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 87.2438 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 6.83936 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 33.0431 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.0353598 LAYER VIA45 ;
  END Uart_clk
  PIN rst_n 
    ANTENNAPARTIALMETALAREA 1.467 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.05627 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.206 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.99326 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL5 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA56 ;
    ANTENNAPARTIALMETALAREA 14.9 LAYER METAL6 ;
    ANTENNAPARTIALMETALSIDEAREA 71.8614 LAYER METAL6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL6 ; 
    ANTENNAMAXAREACAR 559.512 LAYER METAL6 ;
    ANTENNAMAXSIDEAREACAR 2705.84 LAYER METAL6 ;
    ANTENNAMAXCUTCAR 3.38649 LAYER VIA67 ;
  END rst_n
  PIN rx_in 
    ANTENNAPARTIALMETALAREA 18.291 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 87.9797 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.687 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.1169 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0598 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 49.8712 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 245.365 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 1.81104 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL4 ;
    ANTENNAGATEAREA 0.0598 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 52.296 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 260.246 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 2.41472 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 2.682 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 13.0928 LAYER METAL5 ;
    ANTENNAGATEAREA 0.2652 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 62.4091 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 309.615 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.41472 LAYER VIA56 ;
  END rx_in
  PIN SE 
    ANTENNAPARTIALMETALAREA 0.565 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.71765 LAYER METAL2 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1755 LAYER METAL2 ; 
    ANTENNAMAXAREACAR 9.43761 LAYER METAL2 ;
    ANTENNAMAXSIDEAREACAR 43.0496 LAYER METAL2 ;
    ANTENNAMAXCUTCAR 0.205698 LAYER VIA23 ;
  END SE
  PIN TESTMODE 
    ANTENNAPARTIALMETALAREA 0.287 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.38047 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.288 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.38768 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0871 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 17.9036 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 89.5299 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.828932 LAYER VIA34 ;
  END TESTMODE
  PIN SCAN_CLK 
    ANTENNAPARTIALMETALAREA 0.419 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.01539 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 4.568 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 22.1645 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 1.6784 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 8.15603 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.0235732 LAYER VIA34 ;
  END SCAN_CLK
  PIN SCAN_RST 
    ANTENNAPARTIALMETALAREA 0.141 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.67821 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.377 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.00577 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 14.244 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 68.706 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 9.57 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 46.2241 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1599 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 112.758 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 547.924 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.25766 LAYER VIA56 ;
  END SCAN_RST
  PIN tx_out 
    ANTENNAPARTIALMETALAREA 3.966 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.0765 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 3.987 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 19.3699 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 1.431 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 12.932 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 62.3953 LAYER METAL5 ;
  END tx_out
  PIN stop_error 
    ANTENNADIFFAREA 4.19 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 2.138 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.4762 LAYER METAL3 ;
  END stop_error
  PIN parity_error 
    ANTENNAPARTIALMETALAREA 1.569 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.73929 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 21.624 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 104.204 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 1.431 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 36.688 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 176.854 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1976 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 278.737 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 1358.41 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.59741 LAYER VIA56 ;
  END parity_error
  PIN start_glitch 
    ANTENNAPARTIALMETALAREA 1.588 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.63828 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 28.091 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 135.31 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA45 ;
    ANTENNADIFFAREA 1.806 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 35.236 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 169.678 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3328 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 136.581 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 659.285 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 0.783666 LAYER VIA56 ;
  END start_glitch
END system_TOP

END LIBRARY
